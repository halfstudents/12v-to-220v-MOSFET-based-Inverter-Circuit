PK   R��T�FT�G  �)     cirkitFile.json�ZKo�6�+��2��˷n�C����%R�PEr%*�m��^��ؖe9�)l�	Erf8���#�g�揲�Ӫ�񣬛�*��fΚ��?E3g�������o���ڮ���nZ=l�R�*��K)<�z�]&u���0a�2�eA���ݹɒgQ�#��\F}䆡�4B�zI ���ɫ�՚��fl���h&6���"�0�4H��en�P�FaDp�dAd�mf�y�ۆf��l�0�c3t�y͆�a�y,Ά�a�y,Ά�a�y,��4CVYL��X��KjZUmYR��y����|�2�!b!�t�H�rl!�vR2���¶+B�s^�i9�l�ii�l�i�_��i�^��i�]��i*��,���Q\I��*e�j^X&��2�:����Ĳ��w��^�4��i�Ĳ�ri�X�����U����B��Z6���λ�R�fw6�S���ɉ͆�m��͆���l6�G
�)e]�b��գ/�9j����q�����h�π�E~B��*@�ע��='ٷ�l�*������+��a���D�H6�q6:g'67�;cncf�1�1�Θ�Ř��Ř��ŘŖ(�s���V-��t5�\U   j��Ow�c��d=���mz���R*�<��c�jufGކ0��F��sCZ�8�Q�a�Y]g۱�a���շ�_�Vp<)x"@���R} mC�u]x�Ev]d�Ew]t��v]�/�8�%I�w}�M�*.�FuYʸ@"��Dz��y.�����(˼�Q�4&�u+�/2S����B�������m]md�r	UnI�&W��;��<���v�g�9A���2!67��8!�d��!�.<�&�_<�%TF�N�k��e��cT!gNU��h���i7�Q��i!w˸sI̽���s�m�w�{��Go�}����%AO��V����jE^}{}a��9��]��;�~�K��F�yy��Z�hC��y�E-L	��-s\G�լ��/�Z���x�H����[��I!��j�O�OG��JGG���m�S�ֲ���x���_��6WnJ���{�� u ��m�"��dF"<g�ш#0�$	.Au�ǹ�sC`G� =E��6k�@F�p  ���(�i��U�8�G��� �H<�k�>��~��cg0�����za�.��]�Km�3��<u��0IG���A�<M�~���QP媶]֨j=��	f>�ծ.WCfPF��<�B�$:W���Z��kI�?�Q����3�����Z�O�2{[K�~|���_p� ��y�t�aKg�|}I�tfK�V�V�yy#����T'L��(3rՉ����)M��~�κM��ꖫu'�y�\:��}�n��kW�x����~���U����+F�?j�Gu)i��e�h0���}�3%0�t���M
<0z�=�������Q`F����ٔ� F�0;tLb
�wX�^`t���>A�Gs�}�X���z�2�x��O]�Q���D�d8
'�j9�U��c8l�$to���S�4)8�#���·s0�,�D�t�yp ΋�K��+Y���I��K�5�����k��T=�(��,��,r^�PK   Ǵ�T��v�({  �  /   images/44c8d6ed-f4a1-42f0-8f26-136091f6581e.pngd�u\�Q�J�04CK3C( %H���0 (�t#�ݝ*�!H��(��%�p�s�������w��W=�Z�WW��æ�FAA�S��j����PPP���ԃ�zz���;�l�4&���c�*��,#eF���s�I�z8��*z@��$#`&�
���� E�D���L_�W�k���	�;�^"�ʚ�p���,*-++�8�8��75uJ*��B��R�B ψN/џ?ӟ>��!a�U��	��673Lcr���\h�ȕ�>?!��zO�	�����؇\9�P��2�����gȕrZ��?�-e����=A�O�\�z-���_�P��c�׿��F�x�y����J���������_'����-t��pể�p��yHr�y�US��<m���1���KO/�����N�A���]���ި�C���-������ħ�����U>tX�w��.8tM��Ws�wr���^=�����lD��ß���b·���*^|{��h>����X����E��RF��
���v ś`Z�ݱ[Za�u��O*���7��ՠ΋:uf8�͡��Ì�ۆH��E\ه_|���%z�3��c�'������}.Z�|�:�pS}��ן#92n.e���/GCŴEN�!�\2���^�=$,�#�J���Ag���ݼo�8Ͻs�7��8Z���뵮��<��>p�M>�S�N6������~s0tuw�;�&.8J�?v�,Q+r����p�c�m��ld�v�(O~'j*�_�u<�q�7Tt,�*�990��2%�	��n���E�|8h��4��P�%Q5����\����_�*1Zw
3�FDN���ʱ8�o� Q�I��؄�"�?���5�1���:t�+|D�Ϯv���w��(��/N�}8/�yT$��2����jķ���s���T���Q�8���w�Z���������sE��KI�%�4[i��-�Á��_ �6Dt	�����K}cz��l��O��n����z���ݮ^���_��0��0����㬀�4ꩧ<�y4����XAWU�ɣ$� ��9���hX��WZk�l-X��6tdS����%��E8����R T�1�n;�s�i0��<GUl0w��O��0�1��+���d���T�;��8N�Q0g>#%z��D���-ߣ��m|� ~�t�S<��O���l��^���1	�Q��@vv�Ԥ֟8�9���/�K��e���qT�����V��u��	V؍�Y���3h�v&8��R�%�#.
w:�C�\�l]]�T4kBY �� �<#%4�� ��7.ߜTd{�x��V�sX�{��2W��Ɨ��.]�b�ze{ί����r��hM�k���d��*-���,1xn���mq��;$����G��Xy��pd�>�Ϙ�ւy�OL�ܖ1c��ZH�T~s���� ������8�
��ֽb�>y6����r�lo�J0KE�3�}�2c_u�h��<er�Ӧ��)7�����j�'�9��b�H��d����F�ǯ�YZS\�&�t۴_�D|��b�n^GA�4wS�T~�'�TV���9�n-����ܫh��bG�p���(��{�`��ͫ��+��WX�+����ɓ��_��{�C+���� x��_
�_���u�zT�ƈL)�V�Mz跫|�gt����\u��R�X�1�	s��8�R��K/mH}�r�~A�ǰ<<s�-)r$:���������2�4�f�LK�X~�H]����;�/c��ִx�����b]�T/BBw��?�{HWOҗ(�⺾-J����|�U�\9:$F�%��+��� ���%Ǖʰ���R�����,7�<;)�f?��Z��w^0v�xk;���!�l�����+Ij��<<�̂�>>g�=���2m�E�s�h����q�)ؑv������++�0��fC�C�l���֣����4
��)�6�����rn����V�ӭ��5�q��6����*�3�K:�4;����}�������,8T�ի����z6���Nn�%��t.�����5���:9�[KTt'2O�9�.2�F�k�5/�V�7Һ@|��c�� s�V�%K��[�_k��U@'�f�k�t��O�ӯ�6���8t�"xqy�'�S����{V�]H�kyb�~�������o��Ș�1t�`]�:L��,d棉X>��8��0R���K��ѩ���˷�M��d
���ө��Ŷ��I:>a�$��ܜ��"�zIy�]���j^;X
%���Es�q܃���^��י5�MI��LtܟWMx�]�^.D�"
$���5j�ɷ�ac�pw����D��ۭl7U�3���?�t��D�����K��M��³� �D}����y� 2�S�����g�x:�f=��l��Z��el���_��>��p6�s	�0��i���|�&R"٫���}�"v�:o]�����	�c�ȟ�9�&�""�b�����=�7��y�� [:�窐��1�G��[c#���N,���Z��4&z�Ve'_ٓ6x�ص&du�]�f0�O�'�]y���)�D��Q��~]��p�k���H�+�;���h��xFi���ly�<�d�o��L�_h��
�e���X���w�ӄ��'�W{QkuHL��"gRY��y-�W���-.�N������HǮ��V{��վ�
;�B�3�+��DP��>�~�%�ܥ�6�o�ʫ���[H��x+�udж�sU�V�G�Euj7s�ds[N������4�$Kfl6�%X�1J.7d��,�$��go�2�
�M"��c�I�а��Y�zͦmrz� ,��e["+��%8�΋��UZp������֪�Rb�y�Tg��P��ۂ-_���re�Fr}U{�Wm+xv����T�+��>��r�䆋��f�?n�m�H��J�A�6^j�ص�5kXte#3rcd�-�+��y�{Q�E2c��+{Go��gZpf6<[�������l����ܿ<N�?���aE��ok@K�ԇ��y=�iscm	�!S��Lc���|*���y��O5���k��99׿n��Y$r/�$�[}��@����6���)�H����v&�n�c��]0ij�P���<7�x�7��r=.���u�9�q�d7���r�N�6{�b�}1��糐���zB��!���"yS�xԖ��D�[T�1�N�M���J
l%�,6r%�.Z}�<�MJ��]g�ܪ�.�Z;�e�(�b��p���|�d�f5t��xi�t��,�j�\��|��Ri�=���`K�)�D��Kf!ŧ�:i���yXp��à�x����w�H�w�"��^gn�n���y�#��/G�O��63#�|N3{P1�ս�!t�"�{:"3�?5}��y��(��?�N�������D�g)Q�J-a��U�x��')����ݬ�[|�0H�����P2�֋ʖִo���r�͂mV�׊��IT�/\�����O?)*�z[6\�T[�&�]v�Bs��Ju�z�i+�o�.�8E�i�0�{�Ls��4��4�<���XĘGY�;B÷�.����N�
,�2��ղ.>�6s�xۖ�Bt�jn���+M��%}��T��Fa��&���-����޼)��,V�FrJ�(��O��p+O�<?x�S�(wI���0��p�c�|j���{4���ż���ȰP��^� LP���ۆuo+����8�2M�Gh�
U�߰~��ֻ�-���X���:K��5�Yo�S����J��B,��fW{���=��=��=��?&�	�K��_b��y�)nE�]fw?r�M%��/���w���ͻ�6~�n�ɛ����~�;�:ly�'W��Wq�HB}Z�������� %�Hx�/��C$�x�'㓹ABaѶ�X�5Y��<�bA�枙2���������7��l"�b��j��C���*w	�d�0�N78}g �<�N����k/��s�=0��8V�=����\YOd�L���GgD������)2hu�����d��U)Ä�]���*<����6z�� � nx+1{��8"./�AS,.��E>�9:��miCi��,g�ǥ��}o�L��z;�٫�ӌb(�u��ׁ������F��S��6�C�ԥ���ܱ�&6ѷ��b����jyj�������a���P�Smt�����)�rD��eh)Cr<'MO��y/������0V�iC�l���'Ԇx�uE��H���K�2�>��R���N߈g����~*�Qa<S�r�gg�{&�C\)N���0��R���(���W�$n���5YGj(s�㎴��4���{��v�Bl��D�}�2sy�	n�L_�&_Հ���䕵ɍ�b�6�9���UE�	�¡���2�󅥉f�gB��&>�(����h2l� �#���N��w���~���Ȥ6<e�=ܞ�;R��7��N��RG�,4V�7ևL��vK|Į�TT�-�V�njn��T�5Cz|� �Jx+,m*�SVW|>Ř���S��bzSɫ�>|V��A(�-�M�"�#|�i�t��>�4FvIv�,tS��ؙ�i���?�dߏѝR�v���\*4�۳�c�ĥI�E���}֑�&N���nL�<��|��:*p�T��bV�.�W��Ƣ�C�;���R��'jr�J��'�x2����)�90�	 u��+�7x��SB��,��HF
�2j���}N ��[�~�����[5��>W�����\�4���
/v}zک&�f\j���o�Rj��wi��T�
���
�G+v�\���#�ų6�u��r�Y�~��N>..���%ŢK�"f���.N�B۾w3�Oq'Kh=��2�R�G�*o�EX���Pd���0	M�x{6���rq�4��`X��6�(K�<�2��m��.A����
}:$*������>�ɐ�*����
���v��?1�ľ9��1v]�ɬ{ypۀ�����w4�O�,M%�Vܳ%��n�NyH�]��hJf�h��mc�-�t!�z_���ǒg;���w����#�-0R��
	&��Y�1����7e���?:>��\��$�a�h��$�7�O)��X�~mGR^����İ��"�ɇ�p��ՌYz�S#z^{q�;H)*V�׻���9ۖ}�5�>U�)�"��2.�7�}���#z�?�O����Z�@��߁�9Y;gW)��AR�5���yʪ����wR�(�0D����^�p�� �������0t�n�P�;fì+�y$5E?��tL'}~�I0��L��nJ�x��,��j������6J����X��<��YK��\f����T�st/�M K���/�v�MuoS&������z�)�.���Pc��~���T��xr8����f��oߓ�}�������ڥ'�����3\dM`�v�����<?����8FҒB�N�u��R�U�]_,�v31�vJ�'��D�o����o8�쯖�No�<��@@
k(�.?�r�^)���&AHq׃��Q���e�tz�8D��ir������":@��.�ǚ�}�!�Jroh�@���Z�㢛��ŒH?�Wfw�_�/�,]�G*���u1k�\"al��;�5T5`��G���*���o�ϭ���J�:�dT+�ϲ����� �7���A"�8��:��!Q��j�VG�ִ�k�:����.���O�+Hg4����8��o�~'M3���^�>W:Ok���m�J�̾��->��{���X�bN_U"��-�K�n3@]�<CL�f�?��^Ƹ��o	/�g�ο�	\��G(�݁�O"lT�yz�-/[Zٷ��;��b���mNY��lȠ#aB��&�Dg�˸�Fm%[�Sǡ�`r@I
��e{F�޳�7:�z��w�{1�s� �@Ra_��Y"����X����Z@�Q�Ld%P�Z�����@�|T���7g���b�,��!�qW
ɷO
��r\����E��HC��Z~{]��[?�q�/�ުՑ��[Z�E���F,S;�!�U"�d�j0����N��U��?������j�S;D�1��K(LڑM�����F���%0�o>v7jW�4v�'{�_f���'��N\|��H���ji�����t���d0��]�
�,��v�k�ڄ
�a���~	ٶ�x'�G{������N���K�5�YC�dm3$'읰�P)����f�r��7��P�	��|�Ц~������!��F3��y&b ��\�A-V�/l>xg^��p�Y�j-�H��ZJ�]aw�
p�X�q7
�A��b�O�N�dɺ�#;��Χ�c�E?��y\L0�|[4�I��U��z�㨿��ֹ>'h�E8�G��7���X�ݦ{Y� ?�p�d֑4���ǆ��!!(I5Is	yZ��A�Z����Cl���1ր��NKn�3MQ=�TkG��7|5�Bnu �ռ�a=>��s�oX������p�WIy.�z�G����_X��	�O��f�j"���	�z���L����l��M�ϣ]���YZ�2*"9�̗gI)�7�>&�$�����U��x1�	�G�-}1��h�Ld;�\�Y�yٵ�/^�
-��?��������Hŉ��ͦɺ�ͬ1@��(�*Ս�Rn[`Ǜ�Y�N'r.���H�v¸����|��O0������ɲ�zC����ɞ�_獍�A%�,�?DnO�d#r�w�IBoξ�����qzRAV^;��yK�?�'!���k��G�3
���7|�\DH��ŧYkh#��]�6��� J�9Zs�oa�^p~�#�ؙZ��(Y�re��ru�YJ7P5�m�qH�&���wqZ�1� ��cptc�[�gF4f��{�Z��)���/��=)K�q�-��m�7X�!�?4)؃Rt��x��ȬUc�;�ٟ��uԅ�E�� �U��P��Q=Mf���9���|m����_pΡ�Fx�@)� ��W����k��S��LuX�	v���+BK��[�W�3���KV���ᐭ����\���t�W�3��2P��8�NIH ��yo�|Q3|�|Ϊ��R�����F�K�ƽ�"�nς���8�oL����h:RW.�l����F�T�Bhq���s|%�|��=�=]6�Lv`�_XP�ƒ۲����m�M��4��L�@4i �U�\�*]m��P���wn�����o�o�;�^��O ߧ��)�)V�^�����Ir3�¦�����}n�B��6��M�+vm��e�5��Uk��u�O�_
���&}��ތ5��A�>��(CF�����z`)�jDO��X��N/7A�y�����h��,�H�Z��դ���H�k����X4�5�%�o�pB\��X��Z'�C\�o��45�I��]����k�7�����-�|�2��2�qJ���ހ�vq���Z>�X��?} � J��.m�3t��&%(]�������`<�r��0<�(�Ϯ@yR`
�}+�U��Sg�QiO%����	'3lMfx'�L���u���l%�|��z+�m��뤞�]-b羿Ԇ��FH�i֓Ȥ-�9����y��wR�`����Ǐ��//�N�2��*?��i��H~��榽��;�#G��x�B�1T3���x���fo��2�5[i ���Hi �DAc��癀�e������W#��d<.����L�gINLj{�h�~*�ʦm�Ǿ�&0႒�G�/)��
��G/v���R�L����x��U/� ���M�[W��^~�8������,�Q��_I8�@���a�a��{�M��P�9�T�g��i����N�r��b�s^8�_m�v�_�}���`r���w*��AiR��
�ܧ�IZ�O"�}kh۷����*��!������F{��ҕG��T�M�E����V+h��x���c�	�Q�
����W�!�R��f�Ws��r/�ܮ]��P��t^�z���h�8��a��˷��/��=w
Xr���6~qs�����\p�}ˏ}�f���H�ۺo[8��L��}�@j[��K2��������ႈ��G����4��d3��M"�xlr��+�5�y)'�K���f���%�,�GK�@���2��q����f���J)0�1��i�?�"r�S(m���?�M�E��r<�	Y���l�&�����~�D�0����[�?؋�Q�psI�����0�r�ZhN�@� Ҡ~Er��A�r���Bmk+SU>�:����Z���FLˣB=��f�k�� �j1�U����i)��\����6�Я�L�����q���i�I6��G�h�D����?-��`�2|��X�����B�5�LM�xp����?g����g��"qXdt������|S�P�&���Y'&�$\��M"��+&��~���T!�_�e�[����K������2k:e�9×�B���3���?	���Bb���+�H���Gڇ��{��h����P�;�.��T�W�uYv3��΂�w+�;�~
���ǌ��	���ӣ/="`�(DAc�%�f����ɣ��Z�C���ş�'eɷ��M�& vU$�T�P@�]�5���N�D���V�W�r��8ǤB�I��x��rq=�!�{2��O���頌�Dv�
6;���@�=u���H����P9�ߜ$WQ \i@h$I��cy��n:�Em?x���7���f�8dBHxY��V�= q�rм��DD���F��߫�D��F�;Q+�f_|��--�t�{���	�u�󥧌�Q�C;��K�-��%��ڹ�a]���w�z�Y�#}����%�r֕�8�\�v[J�O"�2d��w �����'�	0��	FF ���ؼӈ�i;�`��W��i��4��ۥ����f�F�r�a���o� efmS�w�����L��|ok����CE6�+G��nI������߄%��OC��Q%$����_�����$�mWB�W�����V���;O,׾�̙6r[J�O�K�Y��]��V��	\��N�G!�.>:��4v�H�=1��O<�����ƙd���~���?CP�	`�
��j�m��O�$�'(��n\qGE� ��w�HDP���u���i�^�t=2Q�~����������1�GP/#��;�R�`'��+J���e%���}�f��{�im�(�l܅�ߚr(i��f�S���cV�f�ӗ+֦E�����?�^ ګ�?H�dK}�R+�؟O�A�‎q�k�4��5J,���?kO��âɚȼ�u�K����$����š��KT��*VC�Y���v ��X	���A��{���Cu|����A��rao�����aM���OQ�QT	- �)�¨���`��s�����{�<�^���c����\�E������!dX�N��А�2(;�N-P
f��[��Q[���gaV.��Kȁ��1)p��#�����I�e�Ua���~��S��Ԇǡ�z	�V���*�g�ui4����1�'�W�c��*�k�Wz�jh����g��}�q� v�]<��w��%Qb��#$o�]tn��ȗ���"˞�0��J��� u������c�TSqL�jЏ�ŖH���$,�i����9�{/�����s��_gp�柔�vI�Xv�X%��;�VW|�g�Օ�@�<���;U�h��Pn��Q��Ѝ�3Ŋ��+~�s(��i�a_��m� �L��b��Y��Q+	V ��LӪ[��ed�;	���I}�IYO18�RY'��*̾�!:�����1**�zY���`�9�/�~��]O#��(��[�%�Ux�F�SU�]��Pc�� (5�̴�LN I��򄾃���l������(�@i���ps��o�٘�O(���=Ll �_z��h��[C�<��LP��"2�G`\3�*��NV#�&�ٯ��2�<��$E���	�9�$��	df����'Ŭ]D���\p�oz��o[{&�xD�D�D5ߦ��+�Wk�u&��{�1(h�#�e7%��%��4�ķ{e5�chm���\���.qWa͟�#�K�/�_�wR䴔) �%)��c�\
��b�x���u&S*�bńK�f�cfO��櫼6�z���~�
�O:m��B>E_�,#u������3p���y�i�L���w�ks&�J�=����z3ځ�֍b-�s��*����;雘obb�4���|�|�FUd5�y��X��N,�� �nuF4ɭE@(�1<<��7)���ri��a�<R�$��-��?:��b�'��Nv{+�����^�1c���Z�����d.�>����V��?�(������D������O��
*Ɓ��Zlw�S�*ʓ�/#b��,��5��di��r71�ϮΪ���`mF�X���7,v�k���Ʋ���d����!��r�<�d�Gr�i�����)JÑ��o�G�����|�����Q�k)�UE�'ͮ6RG�Y9��.��c����3*9ҿ%���V��"�E�2�4�6�����?�2�<���c�� �H��y�1��"����>Jz /"O3��)8������Wy�q'�ö��t�I�
���z4���w�@LH�Ȅ�Xe��	����Zz��[�(���f���6���尒?�_��D̄"7�B�zYƆYI����.�5�(>T���*^s�K�P�����4�Ҽ�(F�ĵ��Qs���ӓ͏��*����2'���S�<��зX�g�ysӈ��z4,T��,˸��47}��Z����J�/B�a��6ǞsULa\5C�s�Ϫ���w��FS�YD�ҙle�C�m.�c�F�sd�@:F���֮
A�O"[�P@�û�h>}��D�<��{��p�}��75��ܴe��5(����x���:��[�	��:4��i��;AU��q�D!�C֏�컌��`"�Q ӄ����e��]�w/�m�S ޫ�n�_����a'r����sl@Tbv��2*��|,!�!���l~Oa�&��Ox)�O2�o%õ�ȔWy<�'���uR�Ge�ͬ�la�K$p�9�-�5�l��MaK�c(�e�v��Ԩ��pB2LB���q��x2�\�i},�
A"}���aW��,�2@J���(%oS${��Ä
�TqH�RhX��>��>N����>�G�� �7(s�S���<�/{�S?%{�k:X�Sv�|em��9�����q��=�O��Fo�Ad�<�z�?��/6?�*�9 �:�I �Ty��{5T�'P�����lU��o~�����sA�ތ�����v����ĤA�J� N��c��_��oV�� �^�R��-��y#.���_VI]�ŕ9�Kx�(T76��=�vt�D�d�#�e�h�D2W-�
N���ۍ��?�g���0��G���
N��
)���Hgsx���Z\=��w�m4^���B�Ŋ���K��(?v���տl[�	
�H�t?�m�wE�*���w��J��M��>`������F�FF� ��G�&$��������_=D��_O�跂Mȕh{v�(�1`B��v�R���+��͢Ҷ3��]z,�G&�!�	EA��3���P��~��C��*#$9��%��a�2kV�T4,e8��(��N�
��
1�>�����oZi���@eI =�6��\��p!�v�%=�'Z^y1�������r�_�����A�7�K�1�&ʋ#��3�Q[
��ʵ��صk5����Sʍ�K~�}����Oy#�\��2= 3M��	0��z��ľ��9�﮶	�2�:9C�,�a�P.z82�J���Aë��9ڡ���+;�]��
���o���N~v�s�W����h]��a62�La�X0pQA���wdTg	��tU.R�|��ʂ�� [yr���m7�to\���4�����F�v��<�����>���>>4-\�BL�����Qi6=F�hR֡ƛ��-�1�T#ׁi��Q�sT;������2>�Y�"" i� H����G��e�,�y?��}��~,[�0����l�v�+�=�d��:I��/?_��a�$�t�����~�=�O��8��������]!�P����/Ie��u��1�.`��[יO���;�.��`�`���#�aG˽�,�f��|�USDV���H6�L���όd�.cT�h�V�������3A�*����o�R-��S�lh��p>!�ےy��R� �*iz���#����(�����ѧ���l�9�$o:�^|�o�&�+�S�`���Vt<܋,�0���Ռ����&��1�2݁x�|�C�n�ʹ�:P�J@t&�.�����/q2>���ϥ«ں�m����Hv�޼�E`3T���0�?�x�)\���,�.B���uc���FJ�G4��}-En�L�8}(������������b�Ϸ������e1�lv�jB];�p���*i�B��0��o=���G-�N�d~G?
͘>�k�lZ���߸���ٺ��^����&�E��W�V N�q����N�����HX���M�����gw!){Ys��2�ƥ��/I�ZF�@|""2�)���s�
����B� �����HItg���:�T����f��&���3J>#�~W����)����
�׭�i�{w�B�)H�����76R-�Q( �u4>����s�ٚi�+�t�AL�]y��
իT��v�`��O��Yї�>���~4�Qpt:iB��@~�P3Ѐ��4JAPPc����vSR���Z�ˈ��������MpT-���nHo�BD��%7��@HM��_�#�wH^��,�N��Y&B�Տ=�F��o䐛x90C��ؿ(�aܪls$� ������RvP��%c�<usl�^�iE9�)����:��2�:}����g*՞�E/_�%�D�`�E&��	���4v���U4���O����I�L �7J�E;��0�/�j�ȼ���Y>�)9D9AMi��O=��4���r䛃�O��I�yP�)�T�^4���bɊ�(��կ��Tv������C�	�S�G�c���`X��8��i�+r�=��ѭ�N������ŋ�*+��`���ۏ�<�JM�'�v�JB��yի#`�oA1�F��rvDf�q�����QѼ�DԔ�!�rccc�>H���Ҍ�������)ѐ�.��'��H"�<�U��y�RA.
*H^�a�%����_��Ŧ9Y��]�}5<k�/��KH�!�ʲqj��L+�{��I�E ���`�?�$�j�C $V�G�JR 7��@~-T�Ŋ�pӔ(��z����_��0�G��o�8��r9��_e" ����TOi�4�aM��r[��'�k D��)p�ɴ�|N~[��W�RJ�6���� u~F-a]���㇓�e�pD����G:`+4!$"^5M�̹��i�/4��j[ /G,�t#�	� Bq��T-s�X��p���Ȥ2���>�=LC�?����f9�e��@4�R�����k��륿��!aK!oq���[\ٚ�E�v~>�}k�f�,��_�O�Ydw>q�̛k����g��"۝qa�uF�j0i���p8��Y<�*Ai�H}�H�/��a����u�b���BK�BU!��(�t�û��O�Z�	gD�"3�"�w��1�A�[.:��*����S�C-�?�/d��)g�umu�~�JpA��#�퇝g9Z�$����K�.ylU&G^�l�/d#�=�sV�c�R�B�:�Ƚ�[�b�G�C�S�,�^<���Ȁ��u�M���#"~��U�;�� ��F�J}y2�D|^H�\��چ�V�~��K��Ж��c����t��O;���sl���H�@�@Y$�
$�S�\���O�EY�ʉ�z�'��e���>�1�����^���M.ϻ������t8��c�������~�>4�+�a�	���te	�B�L�.��,��E��a�Q���-���S*�R��NF|��vz���\����5��RJ`��|A'+��v[pHWޑ�d�d�hPS����q���|�aV�Y�U[,w�1���CH5�v�7@��m�<P����Me���r9�^�@�%;�̓͘�#���]�FI�6H�� .�Y��:0�+��Sn�⸘V�O�ŋ3ۊ��a�n��K?(q�9{v~��l!<�����w�E��P������4��q~�>�\�^ ݟ�� \{��y�����PWp�K) 玗�	�qE�\���>��	���I5�
�!�QV6oR2��E_ Q�;����'�j�3&�'��4wފgN�Iujo�}�[�����z����6�)Ţ�R��%a�aYʿ	 ���<�u�n�L���>���8c-+O�
��Qot:�'��`���9��b��dT=�V}3���\ߩ�yͯ[��{�(;�V�^�Z����Vd�����LK �x� 3H��e+���d�'�~���5$.��r����<� �c��``�
��Q�O6RMr�Ь��	�y�E�����V�������TQ;h�PE�N�ն�56Q��8>8	���$<��j{�N6{<�N�byb2��	�2w��:�Je��G�|���M�?ۥ��֣pƅ�w�V�!\�@	�ǞW]NX��~��A�Dy�j��Q<�*4��G�*΍t���`�c�G��$��$�E�SU>�Eh��b+fc��٥�Dt^ae�v��/�''^16~y;��Q*��}Վ�-[��\��ʧ��"O:���"�\�����F�'�!������łp�m�ac��g�q�l�����o�z�a'v�:���r|�s�`�aP-�җ�ͦi\���@�ћ핤�Ne*�v )���yі�qA;�Մ�����ϟ1��	o�b��d���G9T���l�	ɵS����"�;/�����qJ,I-��ʴ+���}!t)�|�U�*Ɏhԩ��!�qS5ェ�<e��o5����	�a50�ʘ�/�<����#ѱ|@��գ�>:u1S
�s�˕)�I�Į�02ؗ�nb5�0�3�����p(������f��>OI��8i�@V(�|�Fw�F��nSi <�VbI�j@�P���V�ۢ��j�����Q���d����7��:��,�
K7����,L���c���'����cf�c����1��	g:�6�a
[NX�i�������Fk˘�G�)VJ�:To�E��Z�ڮ_^u���`ߋE75t�+Y��蓮�w$,��ⶁh��a�kV˼���_�b�:��"{�=q���D;e��	�.�
JJٟu�,�+��怑���n0!������o��a�C����U�޵��B��OI�U=o���_"�U/��ex>޸�h���K���M�G�����aOg2P��M><����o1(�d�����:v�>^�$����F�^���a+��Q��ޏ�+u3��ױm���;a�, ?��zydQ[x�1~o�%���,��v;k��
��ڈ�)��t�U>m���R��bT����W�W^��p�ع���%�$P,�S�Wq��d� � _���=�g|Ed?/ߜw���5r�Z}�{��p2�Bn�p=I�&R���������:���ة��2���Ļ��n�x�Ѣ)�W�'9^l�貧��j�ӛ�kٛW���d�1Q$ߥ_ gF�f��p��ak?���~E1�2� @�dj�e����72�[�JlU��R�wK1�W4�9�����	���9��@|�4��l#��;����cÚl�<Wc�^e�9�Ci4��P��g�N�2S
�G��|͠���@�<P:|t*�_Ps	�K��.����WQ�f���Y�,]t�{@������Zrk�-u�j,����d��6m������W<���>��I(�|��f�#O��?t�ӱhtf�wס��4���%ʝ&�\���\���E���j��\XO-����B� 2���N�T����t0ӛ;�o4�A�k�Bu�)�-.�mۇ�:#����[I��o �u����G�����G��+B�ǻeU9���<D��~��u�z��3Md#}e���Ya�Ogez�Y���Ոo�ؼ�CR��9D_P[,���n�5�n�������z�Iry�"�s�}��򕉶:n���tߛ����vlӍ�|]��Ϊ��M<4����	����^��z=�f��l�J!�x�%��A��.��z���0�ʪBJ����/ET�t.����?���"��>�mPK��@l����UY�n�ݾ��c�;�e�h��u���^A��K��dIO���B��q�����j�6�����<�q9�=�(��{��¸b-���@;?�M��3����T@�<[;�5䩦A�2��%;�n)�Pc:	��`�=��=Q3��TB㙌�>�KF杈,��n:L�i#��7a���$���-΋��l���O�:��x�f�޵,�ok\�ר�h�R{s�R���{9�zAx<�A_ڏ����=C��'��fW�G��g�^��ɠ���b�͐��C>B.b0�i���".eZ�k3j�$��x3��~:~�),�lwW��J���Co�X��gS�B)���2��Z����ŷ'cu�O���e�����?$ebw�'O��y�h"T���>��1�5~$�c،I6��:�|�eJo�̸}Ϻ�l)cX"������lA=��#���%V~F4��'�%���/�:��D蟵�h�a�U�y�)V�c��� 쑹�HR5HG����X�Jf\)�W��(\`�����QK�k�����GҸ�ހ�_�z��L�o%�	FП��Ё$�Sqla�Oso��~�=C�0�t�tw�  ��HJKww��9 (�H�H#-!�R�����[{��x�s�����y�~{^��N�}��Y����6�!3&���@׃ݗE��De�/��3�oF}�5�4����k�E햼�[����5���ڪ������*>\Y�Γ6�p��9���0���ƣ�щ�1�6Uxŧ�h�-��֝�\��I��W�7�ĉ����*�	|[��uߟ����uc��w��!6��ڳ���GK����%���ث�R!!JI�
d#/�z�^�C���R��i+�����>�S�U	OH�%T�z.�͍�=��h�l� �W8�����&���$Kmup�n؂n��D���"P�rY�2�~*��9����
�M���
�W���~����V�Ǆ�I@���f(}�a�=���~0G��x�U��Z��7�c�[<�O҇�r�r(i(�TH���Y��G�=u"^���:(-��l�`EH,�����э�� �gp�S��,���7Fўo����3�8��ߞ��qu�um<�0	��ue#��8���0G���Lq�Y�&� �<w�=�Q���N�ai�L���*��/�}B\�F�(�x�:�B�B�Zo�S-��#�3�:>u���Fp����~���+�ҽ�:����>y`�3�:vG��6��r���n&A3{�T�S�ɥa_�^���߭X��ڢo�Y��4L�"��v��A��W+~Gfrã����PuQM�9鞞i���%ڝ �M)���(�Ƭ��t�Y�K���!�J�/��r4cl[���G*uC��]�g��+2�!t�o�~�^e=^�{��`~�kxZ�{���a�� O��_8~�f�+2��X�f��W��H7 �n*����gw�	^WL���t	ky6�v�v�( ��Q�2���Xa�\h��AX�/X�r������̽�o-J�?N|�iVS�w�urPi���42��N�l�W9��f�a+��.����:ӄ`hw��d�&�7����n�F��9f����m�%��s+Q��kl�*L8(�ɫ������Db��ۤqX�n�v���Ql�Sߟ��nP�=,Q����%4֮���9�6�)�e�vz1�h��g�t�7ڨ8��,��~vG
Џley�_٩�>"�{򄕇~w���w9�T�NA�]��OS]�""��+3��è$�"����}� �gt��W4*zu{�GĞ���J�CN6�mR(j������?ǩ,�u���2N����=�>�3s߼I�2?ߵ]?IIW��<x1c`�Y��{AC�`��P����l�o���kɥl�{Sp��g�ht h��ì핶A�T�ɢ}{:R��HQ���O`�%�$����72�כ��5:t�(�|�ℱ���m[�2��q�Шsyϸ��)�ǵ ]�C��ͧ5�3�W���A�XayK�O�{]�zB|�u���w��3k߆�o
ˋ/��A�����P�msC�Ab��ٱ�P��a��{M�������@Ty'�)ly�Z��o�s`���3�H�G>��\�q59���=��|ܾzǥ1%S��ֱ�>���J��}T�Y��'-�`T�>�������M�A�;LZ�ڠ�q=6rA��_�LQ�y�m�
�����y������Zy� �iB`ص���]�?f(���p�����!�C�z����x���Ap�����J<0���uϾ���'�o� ����f��j�ilkg�y�]�7j����fqz��K~U�����M�`Ϻ�`��|ѳQ\4�,�Á��R( /��9|�z��N�;�k��+*�������5�-zjB��\J,a,m@66'bؠ��zo���63��*`D���w�IG�j�R{��ƎZ6��״s����B����	���Z�N|Ur�K��h���1��i��>ǻZ�q�ON�ӱ	 @�az�L�K�)��'�e�{Y������P5�X�3P��A�%����.��<7UEYW���K�z٢Sk<!�+K}n��w��_&T��������;%A�Ј 0�W�b�]Eb�+P���caLLz �ʜ�b��R-d�Z�0O�|�jU�k�rh��GsY1����h� [�e[���Ĩ;2��s�RнVA@�ݤ�s��tp8Bh�e	��|cGPK�'#r� �Q��顢*g����d�Z+�x��������a���`��yt��;Ld�F���N�!vf l�,���e��w�с�GӉ�c@�Jƈ<�:&8�G!(��8�a� @`t�?.�J��x@b"�o�� �k������lD1c\������p�A1�H�5��	�I
����$)؍�*;*��*��ļC�hz`�d��d��?H�c��U��&6�`�F���V�c\>��g:�몿Y��g�>c0�,�x�ӡ���Ȥ�e�!�(5F��3R��B��pĬ��g��YJ 3e�e�H܎�po��#h���_�x�k��N�j��ݷ[��,듸0���
����ޯ��L|��=�$��^�6w�����H�����z-V�o��\]�~t!oJɌ�YfR�s�t�PΗ����IJ��:}őg�e�X��[�R�����>�9/�`���DVY䵻����� j��X�(gl�·4[(��2�7�X����n�]���R���<�U��&�DW�M�v&o �ڀj4 L֛R�S?�mczA׋���m@t��߈� D:�	fJ�]���<AG�Y�A�@|�2��h��a=1 a$j����~#c������:{<��$��Rl�Z��<Q~�� �d(��⌚ς࿂�z( Hj�q�J�A1���0x��ͦ��9�X�t rl����)O�ZS����	 i�J��@���Q�h; 1�y� ���r���
�:�6���)=fc�>}} v���?$s����&�����O�_����d!�b�T��Zi�Lk{SHp���1�?�^g�<r>�$r��v�PzhkRs���X��p׭t#f����g/Y�	9v����D�w4��껻>���|�8�;�c����A������hQ�e������);٤&���*7��-�V�.�v^� �f����v��M6�X�����z��}�oC8<�V�-T�B� wN�xf��i��6�p7��m�'&�<t���>�&N���E
�Vo�x�Pi�Jhl���5�2xw%��r#ۢ�����6��O�zփD)�	��Z��g��^�z��<z�5~}wNėļ+.��J�~��t�M8+��3~�q�Sȇ���T��,*6�� �BF��d��1r���Mi�j�ܯ��26��+7+�֣��uE�8����a���������̲N�u��<��N��L��m/$�2CY�7����&��8�kYS?�-���@��q�hC�r�f��\��r��AH�e���b�nա1��䍫����O�U	-�;��:�q���l14HR?����շ	R<�o=��i#j��ʪ�`�49R�>���S��M�Brn�k�{������q��j4u��{��I��B/��t����c��둯I�p!��7�--Ѝ�rJ���z�`��KCE.%�SтF~D�̴5:�����x�:P���ui�k^x����������#�c�3�������[ �E�F=��A�����{7�
a���}�1�BŽ.�Sl���	��!��Cu�8R0����>K���(
�WulZ��-������%������J]��8���"�6
scuM�?p�2�g4��赚����y����!M@��1�h4kl��g^��`�iF���\��Ghn a�3US��l��j���7'�5���:��m"��z��������>�лcv��ph�v+J��p��L�V����%�>^W��N>Ea������ܚ��Ε�q�"W�;�GP��<K�rJ���m�<���3ڦ�#�Itu@���Ҝs�h�gC&��Y�����m� �����ھ�/�C���k�)��\�4L`�7o�|�:�UnW���%.>�Z�\�7�eC��_�Je�jj@n0�,�Ra �	��!m&��G�+'臲 ~G���4�9>=�i]!�o;ni{e�Ez��gSJ9Lg����k�2�r���,���C�:�P�I�I�(�MԐ����?���U��A��U�m�X�)�ڳ����������1׾u��"-C�4��`elP�!{��!�����ll�V]����Y� �ݑ�&��PvP����^t)�5+�H�Tw�K��F�O,�����Mij��D������V+�d��X����� Ş���"�.K�=Z���ܕ�2y]̦*8�*`��v2���A�}��5��в����!Ɍ�F�={�p�q��q�܁��x���)l]
,Wa��4&5���}!�A�-��c)$j>ATN�"�m��mZܼ^O�9��:dĖ�	�vX�f[(E_��?�?>�poԶ���
���#>tlqf���q3$�Qʈ�C��Z��-Thvh]#l����|tW�WYl�ςs�ܸIZ�_&���NF%Ҥ��������a�5'MB�(�M�D����6z�WD�P��L��z^=0~^��t�nEn�ݕ�di��,���m�����z�A�sy�oJ{�h�s�ՌA� ֏�d���j�9�X]mRwXQ�(����ܻg�ـP�f�?��n�{8����z�� ��1���P��\=����f�H��y��E�oV��j�i��ɓ.���L_ʸ�\� �ֳ&] {z������8��O�e�Pb� J�z��&+ #;{��6ƙY~�P�E�ƺ`:<�����_�>�D_��f����q�hyg���I�_ޣ�{Y��Y�N�sc�Пn�
d��ϲ���fr�=�H�%��<�L�i-R J�
�����|^��M�@�5gr�|�
�F�9��Ǩ�Il�~�
��2(ӭ��*w�` ~���1z㷄h&k��\��J�|'EF�O��X��8{K�/���J���a@�}96�����%q��^�>hVs#����1G�:�����rc�,"]#��`�����Q�m�"�;�S�t�x�*�⁗I��|�ݦ�����Eq��Y�w@HL
h�
f��@,�Ȋ'�8߄��1�Es<�ԗf>m����$�B���qK�M<CH���Ę$�o��x��}��YɄ[E;��R��
�Ĝ\�`J�|�1
`{{d�UC�{�%��h��~�JGP�4b�0?��Հ���OA���؆����¼~����W���lvK>���PQ��\t]���a[[j]�ē�e{Xc��#{�N �@'�r��������@X�&��|X���YÐ ���v[�0�,T\>�Pyp_��.����aC�#��L���"֛�TT!��D�a�Nۙ�-չf*�,�y/zc�/� ������T��z���4rh����8��|�����O�ĲA�b��(vI�AA27�Rw���ʏpdФ�-���ڼ�?>��L�^��>��#*KF�e`�`.N�9�����J�J�"���{$2��g-����k�"���ʹgc� ����J����l��ݚ����u���Y$~�;��
>y���֐į�S�U�[t�`��Oٻ$�/)_CA��r�i-E��o7�쟺�ɐ���v;�@�J����k���dh�B�CͳϢp��R/k�|��W�U҇�����"�8����	0�7�U�m����H/��3	�2�C�d��W��50�-�]3t����ˁ��| hV{Y����v��%�$��QrO�{��T]Ei�W�������r:��6�������j�z�����^�i�� �9[�E�p��^��kd�d���yE�-��|�����ԁ��3��	�Ӧ�*�&ޞ%������_Z7��y5*NE�<Z���ܚ���a�F�G�zU�0q��^����5·���\���?"���~z>��	H�{6��'u�Y,H�$ B}2�TU�=��@�a����r��A�u�;�_E^Gg��ܜ�nu�᫓1n�]/cT������W��\�9qVȡ{ +ƣ`�'m݌=@�<�|�1o��PûE���H�%r܁�1n^��)	��]d�K/�&�8�*��:�0d�'��7�C�r���aq�A;�ld���J��V��̇��.�>�&z ��!i��4�x��\��Ɉ|]Sz��#+ɓa�.�
���*��KC!�A���zL"��	�
������z�"�z@!Ƹ.I���j*$O-s����ۛG����3h��̺�R��'�3�m;�]�qE�Dҋ̟M䤣�N	y�12��DN�?�T��%9��0ַORe ���&�w��#ͅ�. �#� ��iN?G�pH�]�V	��֪U,'�H��۝�)-)	��J�A&��g<lȑ3�l��=c*ef����xdj�j=I渝h,m���b������[q���<ɳ"�Ǟ�0�����w���v��4�k��� }��h=S�~2NR��s6QH� ��L�"P2H��j����}�Iaw������I��G��R\~��͞������؅�?q�����#g���M�!�s@㍖�M,#+=��a2p[�!T��"qT��A��2�>�h�l[B�+v��ƥ3�w����߼�ӆ��Y���Z�TTT��.!���w�ZMt�d$u��p��\�����2� ���0����QNv��D����u�:��!����]�">�h7r�zŶ��wG�������� ���V�۔����P*�̢�
��_�G M�U/�z�ҹ��ȣ�<�$&L�c��@hM��0��/2V�W.��u�Ջ�]������sM�������7 �ȃY㤛��t�_�#���4�|��>D�*YQz�?��A8o%����F�}<���ri��B�;p�P���o��'�:���u���*���|A���?@+
;ҿ��-,{^���ې����}X�˶���-o���X��4�U�7x�)+Y*���r��PA�x�_�W5dݜ9+"�`:�8�3���d�%a��0y�RA�?r]�d�2�1T<q�@��O�
�Q���e�pl�����Q��ֳ�0b&v��;6�`�:`Į���h��bI�<%}�:A�[cSO��Ж���_54��9��چ���	��'3�e�DW*�4��x_���4�q�o�,��c"5S:����-R)����4-Li���HĖ���Z�6�n�`��ą��Ny���<����{����������6��8Tb|G���zџ頭�R��l��X3�2�.�_������<+�2��f)�~��P݁_M�-��Z�~P�rX����C�jy�Z�V�z��ޭ�.���cCl������U���(ql��a��".�"��p(�L4�a��1S�0x���ls:&�tC�:����J@�h��r�S�:\��t�� Z�� �`4������d���U���QCn�t7P�';骇f�������a@C��'����C���!�ʾ�/gk��ɆI\��L��J+ߦ��54΀��T=�Tƌ���?28M)��a�KJ��@���)�?>e��>��Ŋ/�=����)�V��� �7�j�.��P���ۛ�8W��+gg�!���WIm�u�����8a̿��$�8�T>�$]�gQh)�.��q��P��a�8��� ��)� u���BP�Kػ�S�j�7k��<i��n4A(�_�<*���?Rm �3�9��&"X
� 5����)#1�H[�D�X~����R=��&,&�`�o!Q�L�t�i��b�PJo���~�jA��F�?�^�w���=}����^�O���R	�����NBd��"=���oG����q杁7����wG�VC�KXNJ�y��H���I
��ᡖ�òר�<�ҍʄ��~�T���4������jNޜ\X(�Y�g�~c6<+æ^g�ѿi��P�[z0e��Z�>qa"=�0�Oc��� �"��)��M�M�d�!�9�o���%$�S��D�g	}�g�2�y� РB�d���*r��PQ=+hm`lw0�pn΃�ۙ�@�f�]w�&�=q�Ð���y�߮H�T����%�Dlb�� A�Q,#��7@��iZ��ՈV�bU�AE��Vɖ|�٫e�N���z�ge�[,�a�(�������tEBA�9�QpJ��!��e��s��f�\��&&4+� @�.I�����aF�m��:)��s�L�rvzm3�ˢ6C�a6��� �QS*��?�IC�y]��h�L��q�l3�{�_� ��]���=��b�{���?��}��&i�.!3Tԏ��(�Mn��aE��.u r}��d����1�D�"���t;˵��^PeC��|�oC��ZV�G�buP����>�ѩ�n�-���	3|F}ъ5�R�+����4Ic���F�������L�=�Ұ��y��8�`2�~��Y��|���ur���Y�N�2FcÏ~-�?T,2�Vۓ�e1S�ڛ�S��	���1�%B�Vl�iY~|6ȔQ(R�~���W^�iQ�� 'M?�^�S���M����n4��>�<H�H��v��2]^�KÊ�慷ͯ����lq�b�@��/K�T�����L��z���Pe��d��Q=<)	>��[�NP�tD��h#Z�@��a��U5F�]_�:?sς�E��^;�����c��aW����n�D�ӈQ�\�2d����]k��>M����t�ܸ��'y�3/��/��y ttYF�Y(��o�������"�z&�N�����׃�h���FRO],o��u�n����.��c�C�vH�O���:@/����}b�6�&�R�����i|S�I��\f���)�_y�fW� ͕�ݘ���R�;9]&� ������Ӽ�g�ΖϾ�m���W|@���`qFd�}���<��Ԅ/R�`1劍�nY���߹l֔E�Z|x��k򢕉�z��;wj�$zڭS��z夷8�q�aTvj�b{5����3�u�e�<GH��,F�|'����~����6�[w������q.M��aV�B#��vOw�g�����;�Өj>�j���n�=����"����d�Ezlm�6�f��s}����w}�|��Ɛ�=�l�/�?���;NF�J��/4��t�V�"��%��M��H���n#�t���LW������]��Zl�0�+{�L�@�}����#M��^�gE8[G^�x9-�����cd�K�^ۤ{X�P"_u���n~=`��y��sFg���|�x�B�dZ�[��hR�9�f�B�S��A���*�i���w�0�<qjl,~�@a	�1�W��=�0��r̒��5L%:h7h�&��3 ���o��|g��-��Q�s�oBt�e�R�j����F����W��G<K��]�W���k��*���L���u{jXb�y��\oK�������5J=�ߤ��^�#��M��/e�c���8��e!aUA�d��Z�9�p�ςz��s��U�%�6S��u�<�#BM�8pg"~�q�Q���L�+�2ͼ�c��&=v�و8<�o�d��Ԁ�ȩ��*��-�1iZ^ ��U��o���a�.�­�c.�j������w��㩦�4H�4�5%>|��M���f½�p�>�q?_��7�
����t8�t)p���%�}�)6T̃�
'�A?�;����}�C�(:3CQ|�l�}=�QY��rǙB���в&Q�*"ct��允�}� h�EǶ��h��jd*.ZG�jg4{�T����8�0l6�+�i��p��Ê�o2�ǠA2s��������w�����{c�Ζ�n�]y�KR�q��E�|���K�rq���w.�#�����)!�a��?��������e\�b��E@?.�ޯޘ�3�42qn.ثo��5ȃ9��7q�ld�
!���{vN-�\�R��ֹ�At�7��v&?K�آS�~�K�<�N�5����[�L�c-�8�܆�Z_
.3��#F�?`N >�����TM���4�9�� =M7���Cɦ��$3�"��m&�`|��٘��kО�VdtV�[G�/�?y�T��P�֎���G12n��l������!Dʩ�!}X^�vj�ʸ*6$��T���%:Ǿ�串�|�t_�_��2f�vmV�>��X�mg��i/H:���]`��唈�;��r��p�.v�l�=H�ϴ�H�<�j�Q̕�I/d+�ܽ !�(�n�΍����L)ӿ ��x#���L��ddP�pfu�]v#�\�N ���rO���+㣫Um�++�Ö)4������Ҽ�7~TR1f�u�6���p�<w�����MX�[�CGm{u�ϊw��"]�`!m�	h�B��r��!r΢%�U���hoΑ�����i����Ұ��d�\��o�
�i
q�vo@�9��۪�A>1�����sֈ�T��m� Z�S��_˘Y�jx����љۼ]q��-���`�:���go�Y�����=����:y���C݉pj�\UpPM����o;���*2 Ds��[����X�'�������K����+z�����<3_p���ŷw����f@z�w'S�x��j�m�J�p��6��J�|��ج��8B�	���tU��ֺ�����{�?�M���̱��A���H��h����E�P��������r�Wh$'?q6�����@�Y#�zQ�e��'viϒ��+�p�>���O���.v��-��+�R(��p"�[�YUE�#4�%�����p�M}yɾ<?�����V��������a�i�O��ʣ� ����þ�y=7
,�}.!��
�a�|o~����ֆr/�44^�w�g�K�y���R��tX�;x8VvSe����^DǬx��� f\��-�F1a��������7���^��m)��`d��бrL�u��f�m�7D�3_�������~�G�tu��x+�ɽoCèe,c���xr��E>�^���w����\�яhT�#�\����ZI4f�m������0#be��܉�:�?$O}��+ؑv��gF���$O���@����n5s&����x���-/���9����.v��%Rć�Rӥ���=w� ����W\��*&~%�|I�_�ֻ�k]4b]FԦhV O�
q��/��ͬ�g)~/���BzuȽ+$�ւ1��3�ɫ��J7�,+I�$�#�:��'��O���T�>�O���Q�i��[��}��֞<���dx�ms�����d�����ē��6u��V��$��ʗ��!]>��]�R����Ϩ�xrɥ���*�K�#�U����'Z��r]��	�wJ^<~�d6`��o"S2��E��c��oe��vU���Z�Fx�kF�cvs�*ժ"[:Q7?W�����8y.�u^m�y���dtH�ש�zw>%w�w�Ս!������f�5�>����ڶl�a�����	[�jS�[�b݈B�.푒�\���5^,���L[5��=�ʛ�s�9���~�;���&J�(�`�c><4M̹��<��'��|�'qy2&�1�:J�M��W��vnn�:J�4[,zQ�L��3R֓)���ݪA ]䐜f��v3�H��˯+�I�R�>�t�	��8�?��,jWf�O2w.5��\���<A^g�l䜃q�qu�6��5�L1���c�k���z�7ը:c6_|��O�PqtO��{׸�:� ��w�8�,z���D)�#�l��&!9A�֤B�!5���(��B�	��fRJҀBk�P��"5���7�B����%��5(#��x����|oq������.Qa9�5<E�0���"�Q�F��9��$����l���u��}~{q����n{�ve{Uu՘o"u�M��'t��u�.���[��[�	�7c�F%�q'�T�+���	Z��ɤ�D?��v�<�L���)d%>���2sP��hW]�2!�6Q\��[��Y	g���¶�'�m��VX���_E�}��h{6{6B��գZ�0�b�0=��X�.�}�r�7WO�;���S���`9-��uJC���_���L�f����	���<���l��:ig=m<�q����ѱ:�F��Oy|�A��2ڙOo��P�N�_q��B��;}gj|�����?�S9�ǖ�\�#�"_]Ҧp�Ť��P��|x!X������p��J{�B��u��o:�-r������ʣ�n��H�x�m�ߵ�����YdXG2�9V����gja8��E�'���y�g���kj6kG�^p��'�Ylp����pv��Uy��d����H�����P��a'��ض7oї�z�D��괟3וZ��Q�f��'#�b:����v��v9?�8�"�X>�<����"e���[K��J�LU�#�������X��g?�N�?7;Ή=��������ě2Z��z����V���o�
����DR�-�Gi�(�IVj�����2Ba��0�AVZ ��+���`�IKQ��.�dxOqѭv���é��{Y��n�M7Z/bH�v���u�ꥀ���2��Ӆ?�hxw͇�+ޞ�m�+������PRs��k���-�F�V>�u�{�<�����L����R�94珗�	x>��▛E`�.0��{ko��-#���I-7���m�ʬS|��N���t�V�Y(�҄mN�EY}�Ɲ(nB��N�*�h�B
khW����Ҹ�_,Siˊ���>x$YY��K�rJ�G5_*ۭY��6H�-l�>�a��(�Xر�xq�߭�E�V�������S7����q�6�ϯ7�Jh\����~������Y��a�?7�념�P�4x������UhЛ�wm��cK���Q~����,b�֩��˥q�@\��`���"��o�-~�i�U�Irw�*���'��oF���c,�N,+*��*��Q����7N�컥������0�|eM#ؤ�G�DHb����V�acK�_kT��e�v��ߺ^�*�y�8�2�3�'��՟�UX�����n�;�����R������{���[o�j����cC�>�^g�Gp3�ǳت�W��7�}&+a.!�D�rSh�hI��l�8wD�"u�O��Z������i�W	�2�N&F��۳�;�Fd�\��G�R��7�t���" 8�H����{�������w=	��5.��P;yJ���ǫ�͚�o#֔��~��w��� ��dC�`r��<"� �	�U�����C7���N�uZ��`��=9^�5�o�:e�5��|�(=��+sn�1w�A���r���xV�"��'npkYtF©��ǖ�h��(��!��������O�����e����'���"^e#z����P��tR�����{Kֽ��b*wX��Ƚ1x�ߴjypx���dKM	��AfL�L�'�^�'����< ̍�5�CN��e#��|L��F�?n���0f����i�����W�}͵�����Y��y�F�cN�:���+ݯ���T�ۑ�4:gI���o��19��c�{�Y[��z�̽0�R��C�E��q�xi��T�4�n%�����s��_�o7dr���{<p��(f�%:�x�A0�s��'��HprJ��z��*	�r�6ʋ�t��E�b��3*%
7�;po�+���;�鋰�b�h�A�i``�!�To��ؽo��Ϯ ����00O�V/��D�J�G ��n2���*|U���v�e��UQ����k�a�>ߓ���DD�j�n����!�(���n�D5���F<4��h���V��@ċ�OA�ewJ����z��l��/��\l���+���W��A�+�u6��s��Guc�w	/�:�>kP訧V��Fv���ݒY���	{I߳��6���D#�}>��~C�rGTJb@��{�'���������mK����?�:;W��e|� ���@�V���w`F������>�qhߙn,L�7�c��{�۳ծ =�%����ǯ=�I_��G
���ޓ���E�ZLY������zs�[�kC(M�:şnQ#c7`�j��-�xe�5A������g���^�h�O���������+Hh���%��b#���h�t�=��g��T8��ό��y�5�|��q��]Đ�c=��Gau�Ůa�D4v��Û� ��Q#�w��*-�\��S��A!�0ژ��lX���n����a'�'q*���ْoY�֍Ɯ�j" �e�#��9}%:P���0�ZIC�� Y�l���.�����S�\��(�S���C�A����AH�� �T4��d-B�?PK   '��T~D'�K #L /   images/838b34ec-6803-475a-b54a-babfd323e900.png|�eP]�5|p���w׃���p���n�������㺟z�~U35S=5=3ݽ{�U{O�����/   Y(� @� �𐟖u�V���P� �p�o�ذ � � ��"j�Yg�iD�n4�mؼ%�9HF�C��Bxe$,�2�ه�/+��3#)���:5�f5_��N����`T���T�,� Ӥ�x&��Csb�/�Q�z���!��&�����9���K.�zmz��E|n��:^�(�S������gBi~T��*cI(c��A�J�w�D�����F�ʄe�w�<B����I�ũ�g�H����ϓ\��������0*�3}S-��u7q�3�Sw��H�Ɲ}E]�5�������ѧ��Qn�����'�h$%���I�9��~��F�\�V�"?^IS�N���ۈG�.æ��Y |��2(:�,N��z����Jx
)�iN�ge/T'e%�4#�(SI`����GG���+���f�:�G��bX���C����k���L����{y�rC2|#��'�}w��'��+��r	]�E�g ��P�섀�ݺ�{�� ),򜮘:T��g0��ȠA����7���MM� BW�,$1���d�fT�/���F��f[(4*
�~�J���K�H��B�8������t7j�;�-P*�/���$ޜf��4Ӫ'�OcfS���/�Y��'Xa�Х�m�����e��d�͒-�-�ۧ�7�r))'�C�0E�V��}A���8�sJ�7��E���E8O���ms��b��� �]�_�igw`�#��*�D�L�x���i�'�����?	Ҙb����,��PK�d��"��
�FE����{�v���������cB
b.�r:�%x��f��Vo��Wdz:8s;� �� 1��[�:�9�h��5�]L�h�0�,�KjX���eeur,�A8���K�b��8�ҽy��|9!I{����L��ӗ��
ea*�TKL@F�L=���?��*��e�`���6}��rZx�ZӪ¢+�&��FbQ��l��)��2�l�DGR�ݢ3H3�	ۜ �����ȁc�l_���Q��
P�G1�Y>�mەb��*���D�|�$"_zD�U[&e0�n@�.C|\ټг����4/���ؖ{ <L�ўE*#�X$Y�䆡�DkZH���ڼֆw;���&BA7fW��L�Ql�b���\#c�_D<}^��V�a�ݽ�"`�}� ������R�"IGI����j�K��34"N�͚���ы3w~��{�t�=��>b^�sG�9|e�A�� �:�uZ�$�Ƨ���|y.4�В�� �{Un'ǢCrZ}�[VХ���Z�p� �����B,��J2����'��XF����/���k=YQcg_��E�$����ovP��gA���� rP�؛�
�Wd��Ä�1��(9�td(v��)D)�R����{7?�~Vp�I����0�[�
�|�����c�%���-�^�v������[����īk+V��AC4���ۃ'�A.�
�����(mJ}����
�Eݼo#ca-�Ð�ZfDSF��xj��	h2�؉��Y ��3���$V��7����e&�C�e=��_di�3^s�i"�ez�k�	Sb�M��k�cX���2�!������o�}�8�DWA��-� L2�E���l�q&�u��� £���n���)8�!��0��u$u\)j�-x�����f��$�]�����S�a���7��z�i�ֹ�|ko��<�=�7��n0
��E"�E!���N�Ω��ۄ������l��m2PU��,���$���\��/l�F6�7~�B�D�I@D	�����[�ZeD�%�n�Xs�:W�.:��~7��H-k�rR���%RTIi�#ؾZ����������Y��m����A3���}����돐]�����Xߧ8�۞8��5e&��x4�_���C��q8�l��@�B��sg���m+��)�u��[���d�}F�>ǐ������������}�!�<gg�ﭐ�K�rߓ�j�wm�aC�����׷�/3�ӝ�Y,g�=�b�׍�='��c׆��'P� ��k�X�|�ϴ1�0�:�+�26���������rW�a�M��@2ٿ�
>{T�����
A!Q��z�	����J�R&����Ȣ��.�:/�OE-���=�}�fFk�V�;x�AO����}-����o���#�];�`�/π��vDM���r��GU+-Gw#k�U��F�u)V�_�		r@���!�Iq5��3���[�M�~{�����>Xx3@?����$,u�IFú��~m�`f�Em�0����]���v���?Sk�+�[���Z�G���k��Q�7?�dMA2����}?;�|H}��<"m��Z�ӈ���Lb�w���J�Ú��qsq�vP��aH�����N��|��>�E��,Zͼ`��ݐ����ܜ�2#.��Ҍ�,wպsٻv�ӱ��B�X�-Ϟ{�P�9}Vd���J':Ǭ��i���,X1/Q���9�6�k~�ͮ�������b-��р�iO��O�k��6��Z��u�u��U���p9,��$\�y׀�ϛ%-?�Xԏ�����]�BSd~��<��I	�ek���`-�%���8�E^�̪,٨8���nS�����2DCaȱxg�_8����M���������ɽ�%
9����b�D��v�M���g���J�a���䷣�pНX �j�Ob���C�>)|`���i�M+�ٖ$�
�o�_���M�$���P����eY�"�Dn)
���r�s��Mk8"t}��l[�S�a�v!�Hz�|�6���'��-���&#�1����c�V�
;
�'�I馉@��&���M\0C�kKVzmzH�G�J��
n.�U��&�|BE'G�D���JM7Zϊ���v���*��:B� >�u�@����J��W�bD��7���SA�%t�IQP�������T��Q�I]�cg�V�gZ�.�i�V��s��s��G�I�ǿ�)i4e}��j���)����y�8P�F�3(�9�w�ai���M+U ơ9K�|a9;��4�j����w���ƅ����z�%�m�BO�C]y�2��C"e��!�������� z���uK���Ecs6���`� ����J��(�%�±To�̌"�0��&W_:t	�B��rCRG�]L��r�-�%��C�Wg��*�ls���1�^���EIxN��h|ȣ�,���X����/�[M~���g��uNt�oP?�v��^�7���F>�tŜ���7�,0hߎ4kz�z�l
�6DMa��
�B���e\�.��P�����]�q���h=�����Rx�^�]D��7>&0�z�����!�cAm�u���i���%k�{'�%��#�pqqCp5�	.E�q���<@~���42��k�@��^��w��j�����<�h�~��B`�H���M��\��V9�sI:�4�0�������y-]*'��36��9Q0���>x�l���y ,�n�l��!e�M�d�����#���w��p��Uy���'��A/5/����g3���M��M����Qlg��Mãap=��Wzi]����,�W1Y)���㒻G~
d���'Ї�қ~��oA���7*�o�p�;OQl�P��������{���6�;]5�է�lzO�*�Yj���o��}O���a~k��	p�����v⥄8o�� 8F�U�F�#�
PEx�*�M�^��������_��r_��%&�iߝkՑ�@Ƹ��孹����[Qеq�z?݌�3��Ux��	=F55���G
}߫�b{�dJFP�>��v�UQ���
��6er���-��I���X���<(�?����|�B���0�Q��b�V�p+?w�E1/C�LNs)q���{	\M��N��n�R����2+�Ξ��P�٢�cW�z�'ڥ�]o��%��M���>\.�����L)8{_�B����q���]��B̥HPezh����5��/ p�!��=w�]�UU�,�����U��XBMg�k�N��`�����K�q;Cf2)BV��%�\;w��Xp�2�>��τ G��Qy�C����Rc&SMj���$3� �&Y?�[۴h��Q)��������+����?��$��@��1Z_2���-z.��c��w�.��Ap^(X碪z��lbx�N��^0�/���!Z��PBq�r���^j\ē99UjœH_
��;L:�I[ݼe�#���V�[��J�Z�;[@����O��e��apvDPg�R␃�(}O�#MQ|�ϐǆ	]\����l�qG~�.��G���7����<�n��鮇0��a	�U�d߁:/?2�-��wq�)��{�T�P�_��FS9K��}.&�辒��e�vY��L/>x�p�')��3�4�,9s;�#tqǵ��v���<ekQ�o��eԍ_]R}����/��_��:ߙ�¬!���q߫��Q���T����b<�szl�p*����Qli��c������}mq�~>7�x���������,�ܾW�	��K�m+�#�9��?��|�k�C����M�]�>h�����_)���<�1C�����O���q�����y���>�&�҄|��w�
�7�w��EP�����1���!�=euC O}��~��v,:W�q`Q�V�
�j�.�ߗW�]m�9�����do���ЬK�H	m?m�Y�t�y}1�˃W��.+��+GQ�Π�DR=��C�Aև�$)l�M"��
�8&N`;�VA9�_n:��l_�j¡D��6�����O��D׽6_g�T;@`r��e� 
Hf$a��wu9�i��ppɇ�ܹ� _|�f�I�(JW���a���n��8τ���F�p%�_X��֮�bs���8��`N �T�a��S�=m׼]ٮ>8�N5o9~�9Z�O�]��!���En	�
�3�D^չ].|r�Ϛ����{�b'��s'YZ^�k��l���� �����;�[��6��(o�/50�|��殍Y������]��o����r$�*����,bak�\I(��By3O|y��I~���i ��o��#z�}��%U"$M�A��GN:Q��_���Hf�u�������<�� � 6�^��e�)i+H L(%�Nr4��$�%�{1L��AV��¦�Ě�>�.;�Q�a�80�������3x�;&�hvG>����V`�T~/� ��v_\��?]��xmQr��	,v�(��9W��M6��y�H=CAO�ڧT뒬�f=�X�u �R����5�f��^]����Ko����="��z.֭�_�)q�7Oh=>蜼`Z���)��ز5Ⱦ������^N��Q�0�7� �V��������ɩ(�;�29�������;�s?��:�躩h$���[�Z�7JO�Ѐ����|��ud�;]b���i8�P�w#/_^��� �PW*`�)o�`�y,��������:��ÉQc�V�\����r<�N�5?R?���F�V3f����9���k�B��hH_����)7�}+HgS����a�s/q%�&8�Mh����_?�C���|�����C�Ύ�H��~�.0�o-�%F#`���XmW�?�7���N-)�.�e��T�e�f�+Z>&�b�Y\l>��y�ko��;���W���K��
����~��[���N��������C����M4�ab����ň�3�!�R�d��� OZ�_Z�9�kt�R�ί�̭N�M�r��rŋ����\ߗ��u!�KRоa�����.p������۝c�k�n���۳��������-fy�*>�������Qu˶�nX�*���b��!�h�,��DH�_-�Z�TWЭ):�ʅ)/g"~�d[��f:�a�������_֖q��,�N� MZD%����A�WnՖ���e��E//Ԩ�6��$6I�s��zyb.e]/�a�Bm􆄣kE�k]2�5�(��4���s��U�vs+�� @���\'Z1����1��Z�U�����P�Am�u�z�����n��E��h�匍��P.�,i�ꎳ�Oi/E�ʅzG���i��r�Y0�>�qh�p9����J��1���h��^�/�U�yK�Cr�-�d"e�ϔ=�Jm��Y ���n.��lb��;�LԠ�T9�	v���D�g�l9����i#_7[�5��qwEa�?�1#��}�뺳\Y"��	��?��������U�7�)r�M�-�eg����iB������%�F�����&>�K�Ci�a�Φ2.<m�V�895��VM���|+�h�<�R\�Ӂ����$����͗�7�M��QH�3�VpU��}�K����~��(Gb���67Y[g�>�fx$aQO�=#�7ז���(��(�t��������V_�ѩ?(�{�UJ�RH�	?�)ֲbƑ/�6�lk���%��ʄ����8�DLH��kl�md%��l�~���?O,��^lg%�-��t�C	L�m��.3{<�G���9���]���v螴yr���+��?|�q�m�֕�+�/��z�|�@Ҍ&�aV<}'�++���YGA�"��T���F��(�!,ڐ�O�?��^��wp�j�;�^w�`��ir�1,]x��Kh���b�~�C7+�<w�I�Py��j�\M��b���i�Ҽ#Bf�l��`�UҰc��ĉGu/O0���\H��1�?+c���CP��G�c��X#-���q���j.��f�ùi��a�Q_/����-
�����[�d���?�
����Ξ[�)�7�������٠�Ѹ�-A��F꧴oA�壊�}`�0�� ����B�8?�hs
t�Y(��*$uY�%�c��ȅHy�˭}_~=�5��$��5�G��ѡ�/Ƥ=���Oe�[�K��7fc!�0"��=ى��v ���I_�v�9˸��@4�~�G��*����`I�{��eL�o[Qa�K��0ZTeq�#U{:|2�2
��e)���=�>��6䪀s6�f8�á�/Y�:4fX��Z8�9���Gl�W�!vb���ޤ��`@-͛�(i#Q�+$����*��1+L��O�^0,�I�56�b�-����BC��G�D@����!�J�`_Z�C��>��s�]��{5��1�em*�^c��c���t�����_��ˡa2���˃���F_塡����������$��~���K?�Bg��z��W�	Mh4*��ś�
Ȕ&Ɨ�E�����V�동W�W�rѳaaAh jƳ#��P￁#r\y8��G��M��5<�Y	�e�m�!wC!�M�ե��=�9vd<����[���v�-�88KNYhM�����u}�I��~�ew{mk�������F�L&͓t���.6w/d_���:T8�� �SH�
�m��[����d
m�c�k#'�����|R�F��g�\����8�|F�3ﷳ�:���|��<����n��͎b�������R��I,��0'�f�_�ϻ���O���AfL��k��>�/�ڿeN���~��eQ�Ś��E����Zr�W��	p*j��h�~�ش��t�c����o�����-+sԢ���o���(����W�hHܮk��|Ok�фvQ�Bǃ�2�82mBBe�/�fJ!�zK	\tI��vP�y��PIʘ����*��x���z�۶Ғ����g��bS�3	e�����$[I�r::����Ɋ��!{�t8\E�r߭���O��(��Hغ[�}�>��ex��Vl���\
dE�t.�gj�^�?`3 �ѿ�.G�[�g�������'�~���A�=\���tL��7���jz�?��ި��~�>	ĭ��6w&=���_R�K	6�ȶ2�?��@��h�lo�~å�0ᰟ���a� �@>(�Y�yj�N�
ܽJ�{R�47
p�{'��������x�c�RcH�g�.ό:x4���u�`I�ZU�v�
0,0&�O��������*Aj,�'42`�%LWI�RV���K����@���� ��㢖iP�&�3��!�G^�l�F��;Y�(�k���F�5�wh�p���C(��6Cgf�6 X̥���s�a�)(*O�A�²�` �D�/��6�$a�z��}��A���wE�gN��iײ6�/%OP�T�'��\���vܑ���t\ޗeZ�V����R![�� ����}��sdL������0ɚS#&��<\|Vy�I���.�<����e���yJçl�J�����L4 �.�ݪ5��\�c_���v��ƝԇЩg$gc�wҕ�|ϸxa��L��f�V��e�U'HV��0���N;�6W���bH�x\+ ��o^�1�|%Gx����;F);�-0Ш�5��R��J�E��\R�b��/B40Y8� �h�V_�Y��_l��꾓����"j��F1/f���S#PM�Cf�!I�.Q:��t`:"=��X�h�`Z����������@TE$(׎� �Q��T�s��@�����ǖH��g`�	����D��mKW��w�Xq� �_�Κ��i+��9{�	����	X1����Vy:lmI��^�����b�@y� =�C8�t�>�׀5���k%��@�!T���:+T��}�ec;�����¬���tx���_"��?���p�=͵E*㕪�K���3���k�kV���(��Dp�d�͉_1ܽ}�^45�{�zR��s�!����xR9&�	��I�d4���rMK��u�Ӄ���1��D7����	\���a�16�$m&Ӗ��)�=��!i�!�
,�n����p����މ���3��!y,��?rc�V�+ə�_W=���oy;����|�S����J���F�~~W���\��TfKˉ���:4����f�Kתg��c�>.��tYmȪu��U���}� � ѴNx/���/�x��wn�
��U�FA��\�U�Jځ���BH�����������#��"#��j	}pq|H�q���0�o��^�uOLE]>ޕ%�h��7ic��x�H���D6�.�7;h*����ڔ�w�d���D38��6����C�ߞL��KP�K��(�1������=��(ÂU� ���c,肂�	@2$!������My>�Dib����[��\���M�`�l�E*@�a��������>�n��Rr��\�?lE�_��8P�BCWbg;M$�K��i�n��E����wb�Ε��]��5���m�4*r<�V�b�����I�J�sx���xp«�	��M���MO��q!�^z<�����v8º��P��S1{j����y�7���U�oeu@7a�bE��*�7�©@�+�"�[��|��Zc�T�BIY��%}�GH썫F��ZQ�Ұ��{�X6��,�����c6K�1%�p�ߵs�E�^n.�<C�g�ߤ�ϝ}������cq��4.ۍ�m����0�>h���e�������|ąaS�?E�C�	��Ci�vv�C�����` �.q��[��Dq�/�~#�/	3i�*�}�79�%�Y��g9G,TZ��$Y[�,��&Λ�9�Y�����Z͒}��ᜡ<6��ה3��٫��Lj�X�鑃J|�?UqW�=����_L���$�պP�>���ܿzۋ-�=���Gb����Ţ6v�x��Z<���F�a�/�G�O5�n ��� �F�zPM.E[Md��������E�
����,�S1[�n�sD�U�'����H��W�ڂ��zE}C�9s�7��-[Z?�k��ݵW��5�gOH�6�O#u}�+��!�%���7	���X=�-�|/o�^ǎWU8��_��>���<x?���}���Ԟ.���e*S��q���oۓF� >'��0�o��eHxpc���wY��Y.P�����e���=��ĕzJoR�JGh��_��r_fbx �&���Q���*�):[~�����y�>7�j��EOpD:>�����ƣȠ��=q�'�`�9I �|�1/4> �����x|�����t�j2$��fT�͔[�7E��V��S]X���!�y9[(�7EI�4q_������*&��~Umx��8�~�r��;oz�|:�#�7�IQ��WP�
b4��G��Nއd�7���u)ī�>0lY��a�;|Y�9��g�G\&��W��C�},�F|������3�DpDҖ�r`$�<����cAU�2�TS���Xe1�2_@�m���p�E��c���;s�C��o'�Nu&y>�B�?�%��G� {oN���s!�"Y��˟6��#�*��?.�j⓳7L1�9�B��f���jT_�SW�sk��(��ׇ�J�F�����#}~RR6H(G&��H_uL�t�kHZQ�@���q���ጌ#�R�8
w ����__d�Xv��a��jұYʟ�����EG$�P���ȯ\�B?�4��͌h�g]8�,^���;�?`@�cR��@T��[l�{�Biv��X�B��aSg+#M�ĊL�,w_6��m\B8��())���w(�4�H�rla�G��8�Q��(�Z��ۻ.̄��_�4��A9�^M���O;�躪P�%���V���_�n�َ^�{��L��ao��$X�&��٩��ј��)�h���F�9b~��B�������u�rP�E˶Z'��ɨ��(�)z:rM�Ը@��٘�<�_L�}O4Y�5R�������ٓe1.���c�3��@߳i$X�~���?O�}�z�]K�aoB���of�V`ؕ��48fOV�%4�����ll�Ҋ�8A-#-G9(������~�r����d�Cs!�^���Ìy�cQ�^;D�(~�ݺ��yA��Ϊ���3�z��nl�^oB��(Y�P�6gHٞ�6��Kg�cF�
{1�.�����@h�#�fҴ�3�7��{bK���'�d��_�vI)�V
��Q�fWѼ	�m�<n+�bcT��<�f��Đ^�Y�VS^�T�Q
�E�`�;�P��E����R-�9"�3�r�X9c*Q{�d��r|�A���}�N��,٤^H�
���ē<�?�JN �N!��r�z�+���=*.���:K�q��Ֆ*c�&��
���t��$�Kp9��o�Ԃ��:����Es�%����k;zi$��3�c�$��~S��0��a~��B����-�=*G�P����%:�r�*������]
�Mq?'�gL��;4�����bL ���`ͷ*f@�	�rp��_��o֎8?��+���/R��s-ƭ�ѹL���\�^F��n:�Ab}�[1��j���_���B��S�jYJ��[�ϒҵ���Ԩ�W�w92V��G2� �ݽQV
/+y��?�_ݼt������ٍ�;�]�vI�����{�2K�{���ٞ��,)��
��[���1��X䡹~��*�=�8��Câ7�s�(r%��h0��&�}�r��eHȑkե �n7��O���h�*��_�k<S7cW�p��{������Q@${M��vqeY��O�+���V�v��30SAӽ>A@�T��N��J�Q�[�÷�dt�M0��I��=� �h�4,�#;����W~v�`5�墂����xs'@���V4�����6_��uZ��*�W��lw}�����W��>b�ҥ��R�-���t@�0���;�e^܉d�mÆ��0���C��Ch��h�8�Ήn�myZ�����������	k ����B��/�cډ�.����w�2��p�致ܛ���ބ,�9��V���㷁E/w7�(Zu��o#�q��Ȟ��|�̇����5��Z����vV�
5j1!P�SB=�?���T��jxLf���Gظ���*4���:�Sˠ41+�c��$���n �n߹��WP}/y����c��\���-P��q&��\�Gַ�e�mt�BLk�_w��V���NI��k��:��{�ҥ#?�q��=U�}�(=�z��50Z�=\m���Zl3�T�B�+چ^��W�8Kl-~��ﱐ/-���kK6t�JW��@�8��M�@I��*ῠ�>��o˔�L�W
64��Ы���ZH`v�����A����{T�i��mQ=����q����i@j('�KT�r���b"�Ѣh"������ /ħ'$��";�|�7f��N	f��[bH�Q]�F�&҂�����"���~��,�gK>��7��o�ܛin���'IS��K�9|;J:!=�~���y �<	��j�^%��%�Ǌ�O��[N�I"'������"��fJ���[��4!G��!j�|*�P2PK���������.���q]7�# yh1&�V�F�Ua)�褐v37iy8�o?�3���)B=�#��|f��5�]��wC�4�&Je�a6��Ȕ�PZ\\l�j:B���V$�>�����t���u�����19qҜeX�b�ʏ��(����Pv���ԋ�O�_}�\���ޗQ�?L˳��mr�Qx��YE�u_����W��F����_���ZP���=�����D�|V��^t+N����3�Dc�y�B�bq>�ƻsX��ƧS煺��~�P�hzC*z�(Â_�6� �puD�u��b��]���.�Т9xx\�Z����.�IV�Ұ� ���"N�Br�D�4�QVCZ|%��4�iH����^���^��p͉�*v�-koJ�E7O�|�b�_�DC�!��)���76X;%i��M�m�^T LZ�d�$䖿y�L�oM\�v�;Q	��׈���*�-|*<'�CB����bW�U�Ɂ'���s�E��E]*��l5�<4��>�<e�0p����
_V�\�TG�s������R�y���IcC��q_�����!�ҟ�6���[�[��!�b��6ɕ6�m=*}A�G��W�t^��n�Ŋ��+��J��T}�E"=����bo�� 'H���T�AX�^��n�ˢJ&�	L;?y�"�C�����0��m��;:�'��M[�n��<}\�i59�[v?-����%���:�=>F'?�W�}o�rךMW/z�g	y1ÀYi��	��]�3I��NғT�>d��y�Qj�yA3?j�n"�`R��Q��M�˅��,Hop���R�!��S�Hv�t��*�"Kf�[͘���d���-kkj�]Fˡ�.���6gz���xʰ�ޱ�w��/܄-4Q!� [�Sh�=�� ��)ݝ�Ud�p9Ό/ǒd�������7b��]Y�_,����z��UBY���N��OEO��N	 ��`�Mp�eå�aL�tQ��j`XG|�?T�Iq֡O�\�84&�NhFK]iV�w�^��.tߝ6��<�+-�'�
���Cq�<V��*H������$��S���c �PG`�ν�v^{ؚ��CT5�&��m6^n�p�I��O��Y��J����d�����VC�>��>u�בw���,�;,��roH����"ӵ�ꎋ�'�cq^�/�n�A���5����3�CS1��Ə����.f�h<,V�H��EDF�;�������ہ�5s��C͂,
�7�ht8�(?`"���x�>kg�b���	�&��fl��
f�	klz/�?t�'��fָ��Fb���Ps�dS,�۩{�J6�bD���Zki����s�[P@�9��=A �rH�Y�9���
WA���O���,���:�r�o�\(+y0���I/���ZZ�݁�%��8�C�|MW���N ]��9�!ta�܈�<1�����]��b�d��� �e=��d����9��O@�SZ��[�	��`�N��5Z�������t#�:ĩ�t���ڊʊcʮ�줗�x���s���r�-���n���^7?�ȕG�������湦B�cԵ� �[ʹ�6�����ڪKO��b��{�I!�&ֿ}�~�Z�>"[p�N5*U��z��b�,�1R����˄�^Q�3?~a��C2pw���C�z���o6����1B�/H k�4N��|��B�Z�c1�7��|"�	��Ŗb~����F��+�S�A^�/�N�F���D����ٷ�b�l�
�Q��a'i�\����~��+�=ZIU���$Z�2��]�
8+0f��e�g���.�,bVmX/50;q� L���1�(2$Z��I�r뿶��2��Z��E�C0.P��J?v�tKb0<�=\b}��vX��J��j�f(μ\AN���2?��#�LD<h�h״_�.�����[�,�����\�Θ���b�M���B�­���Cɏ.���oj��-I�V�C���J�Au
	rXg�4شM,	�H.f�mZ|� ������@v�i/�����(6���ǋ�I��)��[� ������Z��&�Ίn�o�_}Zz77v��\��Mj�ڶ�������G�v��Kż��G�l�2�K�ӟYZN:�m:)�0?�PΟ��
�k)^K�+�lZ?�T����OH�=C�������Ⱝ;�$s�X���|QC�kiP��9�߲��rx����%�����ji��/�c�m�}��h6����;�c�[=.e�y�'��;��LS1��^	#��u�}T�},|7|�7�B��0�P��n����><��)��.6kn��"h>�/��#n":� �:-"�b�c]�5�!�e�����n���ף�MѪ븃K������o�HՒAcD3b��햵%G8����d��Y%�}rLy��0�K
n(tF��<iW��8U<M�7�?A����&F!K[;�.?��f�W��q;�R ���5]�pg������/��\�qH���Z"�9��2��d[�Si_�����z���Q����ǹ6�e/��&���V.��O��&�0�mokn�O8n��$���'�C��"o�S֞n�kS��s��8��e�����D\УJ(G�v⑭-{fr
�n���f�d����ﵪnj�S�-1���A$���q�Q�gYvר3γS�pӅ"<��;[�ٓ���YzW�����UQRXj2,z�&OW]�4����Y(���W�=���
�E�])�6Z��C��aļ��)���~|�"K�O,{;]�\^���df��gWp�hW�5���W���*�� �2��z���K�	FO]�j�g�KIFl�ζQF��+.�Q� �g��G\��Y�&3G��T$G�N�|	G���ZǧqaB��$ꠅ��g0�~S�A����qd��3ڒ�ey������di:Id�I6��ނ?V�[�C6))f���k`�͏�UN����i���\�taر������b�Lߛ=E=0R���HU��}=!\��H����q��b$�Yj���ohxjVK��
��\��J�!�"R��d��.�;B�F�'��8I�D,8U��a�?�S7X�{I㘌A�dt�J�����ҳL(�` �0_�ѽ�J@����f��"6L�*���:w�{��,���}�	H�'}�i��Zdh��?��Pq����%?��O�$���Ӈҗ=`��t���	�F�XszB�u�IꭾDك�8�Xd2\�ҬRUJ�6�����:v&��s�J�B���+����a��G�(\zb�ȳ�E�j�!;N=�/zx��Q���Z�j�"D�|E�]�V��$�O��B�ya�7�^�2!��/$�5,�vZ�o.���-�\ڝ��"�T� WK_�����s��7g)����1))�F��b�Ymy+��\����!��o���G��/k/��%�O��E��H3uw���ןP�z�a��F�S�2�Qe��A�}��u�m�n+s�/�a[�MĄ���C�S�E�Ӫ�+<$���}�m6�Y��=/��&�k� �1haѨB���!�Ù�`�M��������<�(��Ut��9�}��y��.v�(dw\.{(zxi	˛�7���=?i�{��}�yR�}����jk4,ެ��d��P��a2����V��d>�Ӱ����T&a�Oz�K�B�����9� �Zc-��R?n�����tC\���e�mfj���-���d�C���5}���f��y�?RSt7Y�t~BsD{2�x����߼x���돷����͏��K��9��U5]/'����vz,�ߖ���~��Bo�SKJ���n�%��[��(���o-@$l��[I��\TDz�ܿ�C<�o#�t��S�,�/\�/e{0E�5Z �S���f&�sr�Y������"R)���R}m��11ތE� 8�zZ�˵|)���kk������a{<t��C"̂6���4L��JLt^�'R<��k#WB��	U�j���Ɯ������h���̚ �F�۶m۶mMl��Ķm��Ķ��������]U��tߛ�?����������8��J�F�ջ/�D#���ȕ�N6��g����"ZYL���ifjI�I�	�>a-!�E�V�����S��'�@����i��i���U "+&Y�%I�0;;�������3�I�~��<"B�B���b�mc��k�}�&�m�7:;�&c��E!}��f��`V��=�hǿ=oP�i�o�m����H�oY���p{5��	���9��N����Y!���+Z��z����
�w�'�������u�{��_]n��Ǽ��[,���%|եF�'4Y�,��Sj��g�CwGK֢������j�m�g� N�X$�Cr�g�_ d��f 4�㢾��y9֌���1��I�p��WL6(G������]����_Y���Q��M�pKuR\+[ɶ4�p��I�$�]������z����m%���)�Eg��������������/S�3z��7 u�}��QJ�%��ު�w��" .W)]��ұo�df=\9ĩX�+�6t77�PI�o~U�{��
Ob�%�ᕌ���p�zB���Y�t�[�e�NN[x��2�M������3g���:}V	0��N��#�����VAmD��;�{�m�hEf��~���z�"���[�א��#�E�7�n��v���r���Eǈ��@�ђ��������t%�a��`T��P��K6�+���cX>�r*���<�5�������v�v|��fi� ���J-n�+��6�O�2��GI1��:���!s��	vB�!�ƾ|.��(�Cדe��!p��G�q�,�'iS+��^�Lr_s-�z}�������w�gˎwGqn��b�bF5Ḵzȣ���N����W4|�n ����r7ӂǲ�uҹJ��V�V��x��m���&1�7��뱆�2Ȗe��nLׅ�a~2sv�)���١�?��l|���6̑k�it pa�1����F��d�еL|N�r�bB�b��18�X���-�?]ؙ��6��5�ʹ�D�g a{!���S�d��s����_Zi�Z�S�	lB��h���M	���
�y��I� �,��%*����|����ͮ�\:�� j�v��qk�^�m�{X���_����FiMO�|w���V�bRap�{$ŲNaM� x��I����Z���Vh�Ly��n�Z�u����Wi�G8��e<Vd��O��g�-ү�I9F�X��
�
H1�IR��_���C����M��=�n5{o���z������w}="it���T�x��}S+�e# ��|V����ԑ� >3tY�B���@dph�Ͳ	
��:�"jZ�����G��@"��+#�k�6'�i��?�9��rF�ID�,�
��X �΀�(0��x����<��)h�S�D`
'�}6Y��0��d�,���F��fw9(^<����b���,����6|p�E8��ps��hT��Ρ��~&۲��):�׌T�,��M=�l��}1L�!NR<�~��qA%wE��Y=�9C*=A��~c��~����&alޞ���/�aj|�Mhpfj��o����Y�F`nd��[�Vc�C4�(=/�"-�&u��9++���� �۹������Q��a���"��e���`G�=ݕe>����fL�e�E�7�[�w=��Ep��8�P�f�/P�F�'ST��bQ���[������@�|�*�&��	�b��ϯ����G�#��ްA4�F�r�7�����:o����~��x�LE�W��������S�<�ĈF���2lv(����
�d<�,nv��	v����GH[�?ԗ�,_bF�Q�ns��%��^��~���`�+.���5�n9^Ǫ�;��'o���C@ ���o�g�@?�T�W�~�#/� b��"Nr0�%.cGhGXo�i�x�u8�@F�1���F!�X�k �ظ�z�Jc^ɥ\�B��ط��<UJ�t�/�/D��������n�~���h�|H��,�Bpx�DYczi
�jz�Ui��]����t��ʭ%
��C� TaNi0��恈�������$}[���,E�ǫ�����,�o�b�9�S;_j�-��f2�H��n+~������H�b	��pŦi1p�����%Q�TGP����O��i*@ߠ�����<�/2?m'�ȣ���Qb�h�w`^Nu��Ǌ�A�'��,�c�G�q9ƘAM��%��h���~)�����z���|˟��"���3ç�>d��O�x�7�m��5���Ui��<���V5��R�h�'��&�t_�����]�~+�����w#E�><�����z9����~Q�������Ɛ�O�W���G�'M\,�����&6M��XOg��}z�4ԛ��]'{�Dz�%���K���D�q�5G��qJ_'�I��H�ߞ�>�;�x���8T�-_��������&a��1*-��>�� ���@��k3fəo�ح�~y���s�f^R�*��`�8��V�`�]�Tzh����c��è�x��^j���Ю=.%0�?�6�9���9�����4
PR���|7�ljw�qy�϶S�,~7�|�3#_f}T�&����5:�Oz�~��=���2vo~w����7Sz�����������E9n�$t���wH�e��t8�&wY�����ռ��'�+QS�Vp��P�(��P�1bE����B��x��ĝ�r:�j�=�?}����x+�%�I��i-�D�\�׸n��S�`��*;�Q�3]s�~>o:�MFLi�8�Nû~�o��}��������U����x������=<Aga�3e��)QJ���=T=�{bÒ�Y�zJN$j���Q&�0<��*y��9�������������Q����د�X�st�s����lvc�a��#ϫ���ﻓY]cX�v��=�b#�L�4�0|������zF&NE}U��l�ޛ$(J�A�$�m�G1�ö���??X���ƖwtN��Ǚ�R����� Q�Fw7Z:Ƽ����s㽺bZڀ�\P�D�wWo�s�\���D��g<�.��\�����t�M���Ч�����7B>X�/��ֹ�]��H���:r�M�x0��C(1L�}�����)�4oO�[ϳ�7d�Rawlu�pb�_�`W�-����TM������|s�$u��۽��Uӱ+�jqR@���Ž���}W��v��؝|H,���}GΎ�}�>W�;�T����WH�m���&D��k�ܣ�漍񚺐)��ܟ>�x��w+|%�_�Bo+g'㖖���?�c/	��bw`;�F%�w�5<�p7R���0��_��1�+�m�yx�y�}�u�Mx"ٰ�|�J�ֺ�%F���/��?k:�A������Y�\ۊ@|�~ٿ�^Q��.��}��6�F��|6.pZ��|��uel�~��l�+��AO�����*�|=9��a�!�~HDw��o���������b�BR���)��ܡw�d|b�y�LClp�L��}| A��p���Y��^�'7�p �'\ٿ��,���]>sE�b+ņ+U�Ls��{�y����K=I��q�q��1�4��bs<�������y}���}A�׽�l��!֧�"uΜq%ky�F��V,`p��>G3$�=@�c�&t��O��m�G��c6G@���T[Q��a*�S�T�?j_�����Wi���s����t���t�%~���o���b��X����e�\�\ AC�8�*����bsKvA����ń�"��e����m[)"Q����+���N�R�|�sP� ⤈;_����gC���aki�2ޯet{�W���Z��8�Ć�֟���{/��~_;߯T��{!SX���@����4�i=�K)�#'�̒DGd��2�Sl�'��4�с~�'b�.(�{�>��n��~^<_�'�g��2��J��B��*@ ��=�a�H�Q1k�tW�,�� 3��
'���.�7=FŠ{B�C�(����9�����W��'�;�\N�x��`i��������J�V��H��fCU�-R����H����Ϳ����`��"7���$6=�y���T�S���@މ���t��J���V'Sy$X���(=��Y/C(�9ЈF�����p�fd/�n`�R~�I&!�W��6U�\��#�ib��72 �$��V!���ڑc�7v0Ǹ��gF%���oO����\�OX��9��5������ ��1q=���>w�M�-��bG��X�;ѥ��kN�\~��<	+z>�_ ���g�IU�o���Fgk�ɘ�ҽ��2��Ky�5&�.����!�NH�s@M#����.�Xd`a���[t�sewYaWV�����32�Rs�MMv[hL����"W����ȹ���en�Ť�>6��m�� }SӜ�,ⓒd6���}p�RA"�y
c;��-�I8Y�ߒ�Ia�I�v�p���p-O�w�R�{���-c�7O����~Q���,X5������5������]���$�s��<���@� �#>�1����M��j��&�a�y�KΛ<k~��W)��J?»��B<��FĂ��Ǵs���#{Lˈ��~��t�{��L|ۻ�|���#���J[n`O{(8�+��%(@o��ҫ������je���֟p��<S�Q$K4�n����@S4k�4���f�z�e��?R����S�z���e��	 �|/gG�<nL,�Wj�!i#Q���n-n5��v��D�������4�	��@,ܛ<`H�2<�+I�8��< 2A��칻����{W�{Y�cW�L[Q��ߠ��y<��z��z���!��-�p,:o9I,e./
K��pd��Z���Dfd�C�෯���FP��Y�sҐ�G�>�~4lӥE�:Ά �3P�	~���$V��B���c��eh"�B���$8�<'���$8B�a5���/<��"�p|��p�h�l��&�����������xSCCb�Ո��P�c8z�A�l���j��VjqJ��Y�[��ْ�����U-���ܵ�t��#�����L`^���֢��<�]�����Ni����(��;��{S�n6��^�J�#B3�;�X$[�1]�G6���u�n��`�t-}���+R7���8m�B ���?1<~�ǖ\���b��\T����`&���'�׎z!���:O��z��Xr����a��ni*z��F�߁=�+�H�J4��;�a�|s��9��bUm����m�T1��-G�s�b���8��?;~,��D��yڇ���{�\ N胱���,�ob�1
Z��ĉ�3LD0E56�f������А��B���O�=n}{��G4�c��W�{����.�#�b���7l_��ň��DhBϪ���ؙvP*�*��v��9��.�a?��=���̰*a�f��C/6G�	C�7���'�6����,�_@�mx�$a��U ���`ʢc�o�l8n	�aѼ��P���'~T�-y�'3;�4)Tr�\���p�sY�w���L�{�vNz���'19�&�0�/b�*�H��x�Pum
�,�c�S|�V�M8���?��9���4"Ԍ0�	��1`�'�Epy(���h��sQMi����=�u;ۍ���XfIi������'A��(æ�A����,O��/� ?�g�L�%1B�U�Ł@��ٺo��㬠�.��2�R)i.R��$zR�N���f���=�|��K�ɜ�����������z+�_+��~dO\kX��oU��^�`3Vs2e1��[�Ҧf�~G�(a��l��f�;h �%4`��/b��O�lؽw��@��!�z`PQ/E��~��H8��Ϟs��U�Zq�-��C?���5�m�	��H.�����(�0�}2����'�rP�ՅK$��k1t�t�C���Mѱ)dޣ,R@7���9�q�g[���&��eCA}@�I�_{V~un����E�1;A��'y�,��'��~J�*�f�z�w!�V&՚�^wB�>h�s�*����}�A����T7����z�wo�i��8Ψu��¦�0�0�	e�FnO�����b��P�k�?|3}d��|�)���P��%��;�S�����60�+[	\~�U���~��B��P������gF�'���.=�D$(�Y$��ei=񲭷6Ġh�$�=��1sm���^�'��n�>���Xy}���U/��!A�e��]!��"!no8ߎ����#ÞgpI��qU�%9�A�ށA��/����f>ES!ش5�m|+v�\1m�+�DZ�� e�`�U�U���.�tI��[�(x�,�s�5�&�����w�q��s�(T/+�vp�Ϙ�}z=/�	_B���I�Eh[4[���:D�N����3��;���!��@۫�T��1i;�-�EגcP��M�l�X�fz����1<�dӹ)���jD�J��<1�wE6�E���?L�s�KlGIң��n;u��$�\���z4�`%hCJ^�g�O����=�Υ[�����a���z;�d��sn����\4��A�;�V˿��$8���	y���$�<NS#5�l"��qU����l�Ώ(�f��V���K�ӫ�R��AN�L���=�����6*H�2R:F��9%A<ǟ��y�F�9�H�U|ّ���2:��NQ�?�bw��K����OY�1;}�ߩ-G���qOX����&9�
w�7���E��oW�T ?��Z������|;Hr09v���fW����P�N�1������l�?��D�C���g �J��@%�xԿ��6�e���p��E�ī�!�\ �iF�"��'��Ip�Rf�AHY�}T���^���19ii���s(ã`��!h�ePFk�t�U�wTZ�a&�=|�Ĥ��_
k���l��ݓDb��QMH-6��Wȿ��4/���tM(��.$Zw��+���1�`-��=�J��6��I�1K�#���f��kQ.@������b��/����ft3�%�!���#�jQ�^�dpE�'�|� $p����慥�e-+���m�wU��;h��2�1g��)�3~�D��x�V�W�{]7� ���1���7d�l�(c`�̹o@�["�Cp� �Fi��D�s�j;��jIg�
˃�Zdni�*iO��a��ۀ=���o%^�����/�:T
>��v��^�*:����4ve�� }�������+M��7�R�%��]��>��5.��__���(qf�Zp~��:�1��ѻ\���>@�#���;k&5�P�+�m��vN=��l�+� B����`�p�8L;=%�9�u,|��G����k<%����������0�&�� X�Wg15�/m�EY�����s6��p�j��"��1�S0�pc����:[4��j�f�8��εx�3�"Q����R_v���kfU�~Q�3' ܈ϩ��tz�_�����6=l��Y��25�]�C�iP� �h<m�î���Ӂ˱�p�:n�J.VGDl-<��42�C���U�6B���~{���B&v�J���>�v���ߜ����i�ϯ(�T(�u��$��+'y�{v�8��``�A!��e0��\b�T����Ia$��9�Z�=��	�n^�"RА	a�dZ�;%[i<�O� K��,��<�d�:�ߌvk����*2F���v���*~@�K�(�"���!&�����b\=�}����e���1��?Ϛ��5��r��0� g���. �<7ZS�N�3��1-6^^�pb+S�#A��ﰡ\��ЮN0c4l*]���wۤM���l-��Tl�
��{��J�Қ:/�M�Y�1��T��`�(.���nڥ4`3�sߋC7J��idPVJ�v]�/a�h&���پ�R�e�E"�{������� �H�R�ĸ�����IP�Fl�[�V�?!OI�R-������f���v��5���G.�����@pT���~Ŷ8{[�И垢����_��*թʹv�����Ҍ� �)z	���<X��#H��_шj�a�Y�V�Y���(i�y���a���e�c*A/��g������b��EE,}?�V���¤ J����� Rr�����j�B�5WY���_���[�Ǥ��H�;�te}��r���V��Qhw���7���%$��Wk�2_�J�(2��LX�2��}�u��ةʻR�3�x��Y�Z�Ji�BԒ�+T�z�b#�
��.T�C5�/���s�����vo7J9X��5_����j��я�NQ?#OR�HQm��=T���U\��ӆ�W���,��@��zG<J�U��7��$�i�Y���k�K�d00�_�k#j��,�֐� k�m��؝��E�D��u�w!��ayS���'G�n�H��`&&�)�Տ^����)ۈ2��YJ#�rA� �Q�
ۚ�}+f+�S�?i���� lͤ�]�j�sF���H�i��K����Mh�4����n.�>X��!s��㍮��)E����FQL#q��FԬ���,�L��ݣ�=�%��>��
�y�[��ʀ_L�R=����M�ܭ�Į:�m�@�?f�	���$ ����s/�?S*�������^k&J���&�Q%�7��g��fJ�o^u�Ha�#�-���zK��aK���!o�)ފ4��f4�%�Nw���[��S�L�"�<�Pyo�i��9.x�|73�L-�L�I���+�c��MA��"-�*޻,�m����-�������t���r�1 ���!.�F���z�845�|޻���D�K�U���΍�B�?������3�1������gN>�C���~Ϟ�(����&FWG�Oק�K|dFC�Au�+��JL½iw�۷�L^D��#Ys�V�;p�>�dX6g��+��d���ݴ+u�Z,,x��떽��p#�����߶����πHx�O�f?;D�d\�����j%�\Kp���!�D���r��/�iG!_5�7Y%���aq(�~�F�bb�~�lOz�tB�d��y�-	��f3 e�m+\�H�@�d6KlG�ʹ�}.*�%+�j�Ajhy|�<4�.rH����ϋ_f���U�56+����{��J
S�������L�8c�����/��U��T��:o������\�k���wA#L���zk�6���5������8�O����\��h���s�hߋ/�w��y���LN��_�zڜ��'?3#�ڈY9r��Y���C&Di�麟�2,��7 ����"���_j>�2�!��l�ɴ�7�2��'4��V��=y���&��L����ӱ��~���&�̉��~S���gD���{S�`��֏����~f�z�G�եШ���yZaQ�v���^�r�1�.�Io
6?=���Ҹ�$j����oٲ)ZN��;G�!<�*H��
��4��1���R�FFA��o�K5kX���Z��X�b=��=�aZ����q��:ǭ���\k��g;̊V��*���Dm���5/!�������Y��mh���,��G�S^���`fn�?j:\�m���ϳ�B
���EHZ.�����ɿ��=__�����I^D�e���y>��Qʢ[7���������
��[~��A�}n�֥�+��K�W)�����m���.���
�Lu���?�+�
Đx�|+*\>�A,�O��7ԩ���q�������`=#[��G}�vx�����$k���Xt8/����ſ��9�Ɂ���t��^7����
�3� �tb���j=�G�_CJ���	�~k��!����<��`�-	/���33��?��bQ�S�P����C�i�@dxJ�I0Mn]�}/�W�ӌI@e�x�fC��K���Y��j*%TL��/!Y)Q��"a�J �R�'�ǡP���'�1��{���l2�!5l'
�7��|�+j�y��+G�)/}�E`���v���&<)����|��"��t�̵�hp�z��#s���C�����/��~�,��WIr
�a�Y���?�@�
����#D
��^z����e����3�$�<�]pN�Ȩ��\U�1��B@��*��9_;m�Ƒ�/ ���N�SC�s���0@�[���OGsq�az����J�Z���=k��uSsEuj(�D>��|�iI�ڢ�����+|0.:V%��<ߖ�l�|�r`e��۸QeL��ԡ�Q���X��(Q���gwlv�(,aJ��p~_�71�"�	�SBn�m�kȗׂf�*(�U�¤5�J���m�c�uh��S,0b�,S]���#��-%�Ն-�7���t9��8����e���$�߂R̚��-_9���d�`�\oڤG��a���F6��J
��%��$�`�-�jў��E�{8�i��?(�0���,}�y%zYĔLXa���Su�6���q��-hB$��k�<��э�sƛ��GӫT�ߤ��+s���̬;�����|�ey&�n"�r_Iǅ�'��f���rM��+_�P�--�3�I���Ö�z���k��r�ً�;�stV?C�VJ&[�/�:.����Y�K��,�2��x[.����s��6�\����p����b��g��ꢆ�m� <˴���Yˈ˓���;*4��m� �ZzA�O���=lQ���8�&sdt�����'��~�-V���a7��k;�v2>�2��D�L&hP2h,�����!3.�K�փҵ�b	iLMYY9��5���Ϩڕ�)!�b:�ϸjB�m��F���m�2 =�s�t�=�P��E�U�gK��	�B��Z�T�y�(HNu�+3�����ɭ��8Pk��Y���Nzp}�g�~�Q�i,��6�9	��S�E_nT>\���=X#�LO{��L�:�����z�<�H'��y9wJ����K��~?r8�VBTc��|���0ω�D������),���^#-����sܛ|�g���Q�;��z�9}��1F3!�i]�д/e@d�2;����Ed�Yfs��?����n|/����v'6�,J{9d�v̘����yv�����'�g��.���}�K�>�FW�������g6�3��_D"�
O��GkB��\M|��,����B6����Z�0�CS�Ѕ��~�(��!����k^x6��s�v�m����ސc�]���|Z��|+61VT}�q=�y@�&�a�I���ӡ��v3��W��:P��Kz�é�$�Px�56 u���@���S�N�s���j]}9p�A��c{|/��æ����sȧ�kH�s�
0x�b��pz���e'dVj`���N������AR����F&����S�X[M��~H@$T60����3�#�c7e���.J0�B�Z�7Z��,�?;�O�0�S��Vj���)�Pݰ�$eA��)�3�� �$�7����]�lz��Z1e<J'��j�ީc�j.&&�J�22+���w�bZ�a�ܱl�X�Cg�Gs����L�� ;��Z�t�dO��U��F��h��9k.�k�e��L�F��[V����X���}��r�%�d�o��{��"����|�/A�/��C�h�6��dd�'�b�VO�W�z#-�3	��y<	:D�,�0�{K�|��WpG�]�:���_���h
���=�׶�a��w�v��H�"����/c��,���Cm���)q�c����
`AY��g?�{�r�9�Aڪ�M'��(���
����M��9*u[(C���ޠ���m�	\VjG*�}�9e>��o&����D��Gz�$+�9@	>���6*�|����@|5/��iu�S�Fs�SK}fy���t���01�!�op�JT�����H=̟}S��t���Omu�v;�C�$��1>���@rn�3�"g�9���e*��4ye��R�WV)7�N�.�ǃ���ey�0O}���J�cW�CP����ֿ?�t�v��&���l,�1����6��N���V����a �
U�S���X�g��v<�n�ͭ<oA������,�Z���-2�k���oނ���s�rg�m����>+-�,���ǂ��ֵ���b� Wu;�5�܇��s�(o�m�>�$���9DA���]R�{m[��@R3VE��O�3�g�>��F�H "��x��9֢��[�hP��,�+��b�(4 ��R��fQT�,Z3�U*0
Mޱ4���zo��!��\�;uf�/�p�[oڣ�a'&"#����>�8�4� {�g�1�%O :=�m�M0��`�� �E�`СY���j����n��WiR���>��Nez+�[��"���#FR���z�v0�
�^�bxtz:Aԧj|��U+l/�
�����\�+��^��O���g�b�.:O�}�y����Tx���P��K���3�� �V�p��MЌx�m`�f��S���O��;�� o�۳���%���L�s�FC��3��(�:�a�p�I�=ko%47���O�/�����G�Y=��.�eW��E�ܤm�Ο<n����~Z�i,��䙪ni<�Z�Y3�5&�W�z0U�����6�	^A�O&�o���U��Wη/J�Q��R"m;i4�w�k����LI+�+c?J��iPQ��ьr�Զ�����A��D���/�6kHSx[�D2NS�9��fB��IHF�W��hz�?&�ɢy����а�,�2��UmV�>�nϴ!��Uμ�7��7�m��{.�j6C���cݴְ�^��F�j,ɦ���Z���U���ALꇥ%w�t��]>�33�d���W�n\5�eJv�����<H��j��D�?-pܛwG3�TN��Ƃ�|W����^:$�����o�����`���A5�z�r'zhSl�Q�A��\y�!�4�9e��:HoQ������ iF��C:�t�M����h�Y��"]�h^Ý��^-�ț9���W��So���ȓ\��L����X;۫�<����G��J�
=�����PS{VUC�d��ぼ���d�K�M��w������@xXZԭ��J�RnӿT|{wǗ���b
����1�C��Q�`� `���R%+Sɱ¡:�!�	�A���*�S��a�*�	 �P~�Ǐn8��q���*JMf?��ӕ����,@Q�O�����@UP[B�fl��D�~5������LlŪ>��=�	L~�S�1/	���M=g�;���B�D"��E�E��c�=b'�1�M�^������X���Bd�Y�r��
F����*=9�o��=PW�o��g��9R}Om��D��4��Q�Fc�hhh�T7���a��J϶��s6��فaD�[y�JД�=�)�5�4�U���߂��;k�9޺�]m�Ʌ��x���]�!���?��/F�C-�O���9����j&�@I��ނ�C@���Y��l	��v%�X-v�Px�˄d�8H�!��#Jqwp��nv�`2��A��Ų�&׽�Q���V�3� ��+>�rpk��/4�l��^f�ߨ�]hx�Qk�H?�,�`�G!���Z�F�4ݧ�Y������3�M]h�*��p�)j~�nA^G�9��H�`�,�wY�����I���?@��m���<u���>-ez�:����F�������y"2NWd��	B��\{��o{5a�6c[�k�ʻ(+gN��;.�ݏc
K�$]y�d� )��id�['O�F���/W[����@x�0V�kU����Wz��̤�����NH!����"���(^gS���{�Pm�b�Td߇�����Z|���?�5cր#n����Sm�~�9�e�����:��Utx;P,XtT�M�w��^�2>�� G�Zv&��6��Ǌ��%ǅ�|�|���k[�F��"Q~�j5��m\��q��>I	��◑�wUWډ�����J2��Ս�*���m�M��"��Qq��z=����� �\��<`���C�D��$i�(]�ƂB.t+�p�0��F����$�)�终��KB����C+,�A�]m�d��qg����k�V'L6-���+f�C��!�]�^"&&����(�Q�LF�E{�])Xn08��2� �"`~�vZ�@\g3SS���H叇C�_w���eH)#w)�� d/�ۗ�`�PRw[� �Q1�\�i1Uj�x:���Y�"y���'�f�7�å�]�}+��R~�K��m�ҩL���(]��}lO�n�ؖ�Ed�7G��o>Hb+O4s���������6p�j�$w�d\��XM��,oU�����g�����Q��|�����x�e�@n���^��z��w�%/w�q`Q����0����]W�u6֭�<xhQB�$�sⶕ_}�����!�G�dx�e�or|�.��Y���-�\�	J��
žj@�Дi��d���>��+��D�)�J"r��_�
)ck1�>� �m+��2�L��h��e9k]�B�rm�'
#dH3������vY"�b^,��2�$���yF���~��u���x���L� α��_�������2�1���Ӄ@��o�z;�����Ko�����767x\�+_�E�<�Ӑ7�M&�N�R�<e7�z)'jQJ��W��s)\)�+E�u�㐓
b~f�~����ug��S�x�އ�>��6�t��E�X�7g1�&y�����*r`�=L}Mad���:j܊�s6�aLhR!l�Q�����~����*=��>v���X���$��@>	v�u�u�����VzBӃ�b�e�3gt�h��̧��m�b�M�AMW���J+w�!so-~Z6� �)�P��ddIL'�Z��k��ةI��z=i
aV��-fk2M�`�t�#�w�;����gQ�S���#��Ãp�#�H&Ɔ	��b=PպoY��-�$j�V��k8@��0;j�k�;������_�	�FdU���f�l�_�l�}]jo��F�o���4n���Z+��)烪f�aXM���>�nc,�Ȝ��`�kcJ��Ajٽ�4S����>EET�Ό ��Zu��H�����J~6��Z�Ohަ�"�M����s���ba�0V�wPވY�$�+Κ�+����t܋�S��:6��	�܅_�!*_@����L���{2�:��`ə񘅡64��4�I����t�dYL�)����8U��zjlH�9�!j�r���B}\i	�\����e��4���-6VҤ��8T��L�����+�5�Q��ث'�H�?�!�:����Kd�-b�  B]����n��Mjc)� ��	�r?x����� ���w��x�W�&�i�3:HJNc�t�(
D�6�4�%�J�q���B�9}����k.��l�}T�=�C5��4К��nFXUN9����/tx�k;V��Kֶ��~_�}o�����XT��v|�y��ꬸd{\�\}�ߋۓ)$��[5��X��U��QN4Qj蜺��7%\9�(ih�WK%��Pr�Z�Pk%�i��(f!��O�f�������,��%Oh�
Kx���ƙ���x�~��?p#�GV�ZR��C��U��F�v�=mOeW���\D�J����h���x¸ z�M\5d$�)�w3��؜�H:���f��� ��8c�؆D��Z�i�a.:��tc����H$�s/q�r�/$Gѽ�ΤP�cڤfk�����i�ˣ��i鞔+F����э���> �)�f8��Q�og{	u�]�;��F�*4�kU�~��VpL�� ����:6��]|�V{fYb��Ȏ�|�O��|l8VK�q�����}t����{\��5YO
�a,�%[)}J2�z쁑Գ�޶�+M�%S�pW�u	j���G5L7B��{wq���>I�fU�*��^�)�T/������ of��/��A5��H����^�j��X���Rǰ�+2R2�u5�Cu��hԻ�(���ܴ���|L3�NX�^�',���d}vk����0�"��l�?Ob]�mӄ���������S�_I��W?���]��������d���P��ߤ�}�P#�r�y�v���~ܟ��s�b�h[�[���-�B{ ����t����T�L�ͼ��&�AIe��4��MH���u
��� ������?iH��q�lF��V�ߪ�B(c��
�ɎR�����ؿf�<R���(!��JF���e�e�a�Z��7p=_�C]�z�7�L$RH^m����o�$��Wů�@��f����s>��+�s��z�!�+h ��,E�������Q�����?��E��Ss`����VI��qJ@�����}b���KY��*b���DV3@"��L��M6�<,�9�f2�
��+?���)�G�P�X������ �@q��>��S�%�T��s�?o�gk��B�� �R�C�Z��߅H/�?܂�uX�
�*
��>Y�� t��m˰�p\õgV3xLC�$"��z\���sȮ6.�`,u7�tB����9��wuLX׽Χ�z{��1F8� \�g�q�)��F�c� � ��NNi��8γ���&˹q=��3I�L�ٮ>T<��!���IN�� 2 ����J�\&�q:A �d�0V�m &"Dr;�)ş0� �%��Ձ�J��8^R2�	Z���c��ԮV ��7@6T��8Dz �X��=�$�ޯm���m�ìIFEp��lԠ�9�wz���b���ԇ  z�eE%!&�� d&
p!+������r)�Ԍ�d��!2` p�ʊk���s��xQ�dDt\�b�A�'�9qY�%��%�W#� �\���y��A�`8�ᤳ�AK��Y����U��! V��w�f�>w5��8����&_ܗ��pr��f7U� 0  ²�;����q)�h��=��T1�`Vé��� 	  !E���t�z�:�)��w�2�qlU�d����[��
�U�<����BDaU��=+���,뵡^Z����t�D�%���4H�U���-�`��r~��)&��pgN�Y��ÓÎ��#q�*�# �u/v�U ^�9�麯��v7$�|EDwZ��
�,��&�^:6�5ϮL�Pr��N�onIĴCNTQ`0_(��L��=#9c��� $�����@z��(P94@���[ �-�wsݽ]�6~Z@B 8��4�wE'Z���h�����|�-�������q�(nHľ�w4�X�]K �fꇋS�T��.BHHL
�ZG��+]�u�yܯ��T@�I�� �]�d�%S�Z��t2�r2SȤNe�eװ�0�F �ѩQ��bWm�=�+���~�!;�w([�z]�A �S���N�て�Ȥ,X4��!��jG��+��eΟ�#�r�'����3��*��;�қ�<ѓ;��r��$���Qq:P!��@�WeFOs!|&	�` 0�=�#~O��,H���%44D��lruruKh}<��>%����P&�z'���c�A��&�~��:s�h#D��\ D�mO�*ђ��� !E������5mL$v�(]�rcp4��E�a�pD� ��E�q@���TSx�H��;�Г��N�c� �i�G�ޱ���}�w��� {�1�q�<�f޸��GTc�x,���߸`����4��k�cYY0]��	�ن�Y\>�������3b�s�]G�����}r�C�#�Ѽ�,D~NF��ԓ��k���H��*�4�2Ķ@�&�ƫ\G�C]?���r��0��bs��]fK '0���B��.)�Z�c �Z)+�k�ߵ�G�������be+��g�P�J�yxxx,"��K8#�P�`JL�c��''�:% ��u"����~!B�!�i�mM�{W�6�';��|r	�N}"`N�!1 � X-�rsh|m]pC}��ɵ�D�H�*��3s��񷷭���O|���~ 8�/���/��e�ȟ��j��A��]+jtn�BH�������5��ж�.�2�3:N,g�{SM�=�|��Hə��0!eJ�?�9�3�ZӼ!�*E~f�.`����ߓ�d�h{�z�m�!�qHjr:�����N>Q��%�`7�S]" �;����ڀ�����m�{�����[�[��;�F�u�+����yxx,/D��!_���|�
J��/�F�-?e���Z)�&uF�ki�X7�N��kI��VϜC
*�����/�䫫�ozs��P~�r��<��G�~��ʽ_ٺv���Ͻ���>��#鑕bk���g��Ɍ/g�ܚ3��d3�1�;�ӯzN���v���h��i�'� T��SEv`�z{�o�4SytA�qp��``��ؖ�p��*& �-u��MY�?5^*��\�Z��_��5��8�U�����'a�ҕ B�Wm�	DN��3��B��Z�̢�i��Jxcl��*����sJ���M���`8<�Oy�a�#�+� xx,rhS�뫁��9���(Jd����o)|�8�$�����_��)U���Z�t5��Y��0,&"�E,w���H�`6&�J1�6��կJ'2��cB�.�����j�O��	�있W���!+���� �"*p����8�|��=��L���{�OBI��ݲM�-��B�k�F7�f~2o����� `�Tr�h�9Ӭ=ԹpX�e�����(�T��@���s`�f\7	�u��qKl"br<���p�W%:�M�LP�]��V�p�﹝�D{K�uMS|8�Z�s{4m!E��"" 94�p%�c������j��aA�;뿐1)�ƯE&qW/���-ksBJ�5���W�ݶ*�&>,�sI�@d��F�'u���'5�6�O�g����],��W�>�_��r���&E�'V9^� �R�%09Tz{ �_�-vAց�C�@X��F��-:�\����+I������X���9C��HO;Tl��C  ��f�[x����o��ȼkN���m
��v���g%��#�� �B��[wǆb�'N���aK����c�B.2Mk���z�������D6�?c��že�ƭU���C��tv~lUfu|X�VQ*��>���n�n/Y�`~lf}�Ň�����`���m�m��N-p�5Y�"��ZH�*P�	J�BzA[q:h:	'�{v �(�u!I� ��j�z9����Rh��mL�D�~�6��ur+��[�x8�9߰j�w�����^~�埾�Ӿ�>۵�k���"!��-q#S�P(hjt��e���D�V!UC�67��*t�OK�E�d&�D(0gmb�dwd�����[WEebNܴL۱�>�=7�c۶'�j�!�C�|�X.^e���M��(쩢� @s!r&~1Sf�,��-T�Y�cB��2   H!9��
݈����x����/�x��;?�����M�B�К�5[�n}��G��G���<j��:����"�֣�,�!�BJdsi�G5/�Z5)Q�4���%l�?-&[��������~��w�;�Н%vp�H(Y��{������&x*jQ�����_��㪸�I��暝N@�y(O�W� �)���&""DQ��#��
���^@�StE��)4�r@ώ����@A��5-k����[v��W���o������׽$t��� �߆Xm=?�E��-S�Tu!%0����V��~�'��oz?(��O�jk+f��?���v����y�>'ns���mC Kк�wB&XEE	�ǡ���s��J8���ED&���G`�8 �*W��Ν�����?x��מy�G~�����lol��~���I�����qa�[% �M��xx5!E���D���bC �ȗ�� f7��v4ŎOԏ�%W_�]b8q˱� ��� a�A�:��$�T�]�; Y�/��B��~�1�Q% �uM�� ���F(��jc�5����cN�n��W�	 ��&������}�����{v�������_?4pȳ��� �m厩u�#[�/wu+��\���b���-�H�"�kҸD�Ȭ��䦆��S�R�jRK�j�5ڪJ���%�4�r�ʛ.� (2D���͐�6Uq:�>Va��(  "�1KY#�
�-���so�EHq�`�2pH�ZjΚ�����(�7������-�-��n{`�#�#S�)�yx,DF�63��f�#�oH��4��q\�١*BJarG8��Ό�r�.-�'&"RZ[��Ǉ�S^RQM�����y�w㍅r�ЉC�����\�{�]�H2$6ByO��(��~F�#������I�����HD�6����ae�~�9���~Qw���i�p~�ƕ 8�9z��o<��s�gn���w����E|�����W��.%�qn=�Z��د���|������P�)��Y�L>��1�>�  s���pXA��{`"�>�o|��� hU�h(�����:��]�h�"I�X�}���FO��2�t��� ��M\C ��̛��к*��v�4���|�q`�rh�-/ɼ�U����_��D&>������>�s8ce<���8���䫅S�Z/���ܬs"G���N���˗&���B°_[W�'���D����
@�r���5�r!RK0s�*�X���f/�ׅ:_�?>��ֆ�ʿ �O�ݸ��{��>4T�����^�����6HVSQ>"�al.���a� $v����L�nK �5���
j]��L���\3S�W}�;% �\�HR��t�����`0�������ҦU����2�2�
>�����ȓ�-�Jl�$ N��)}�Wő���� ˶�e~!E����@��֤2b-v�DL
������d'�k�N�ɷ˓���B�� ��wv~��9*_2��+"�"��;Khk��z��lBN��W>蜦\��x�1���-1��y�����Bh��
�^��u��#F�Z���cNV��z� �QP�� @�k��Tix_~�{N��K ������,�'� �rS���h(�kݮ㧏s�́zx,D p������+Z��rhS��5��=hL�ʝ<p�s��B#R1�������/�T`f������o����	K"�n�ţRi����y�d܇n������И5#�%���1�*����d�ǊF�~z~N��=Y��N����/e�αn����v���#\�|Uk�U�_+������F���K��K�� �����)����+:����7�7��%z���   r�v�] ��D@���x���2���`P���U[82U��
uM�;���(K�u�Տ9Ƅ�z��j� 6r�߽8��)�t���v���SN�'ɟ���G�6����>��18e��D9�4\�7��V�C� �9>��� �����W�����n" K���Cu?{/3��S�� +��zܴ������=���H�9�5���`A�.���Ւ�p�9����FMS�D(�rx�ވ�,�vDI	o�B���[�kJ>e�Q��N-[_� p�������o{p{HYd�#1�}�>/��cN�����`�0�8�B��7�3�C�E8 �?�v�F[�$"������J 2@�r�S��+C�C��T���pԂ p�L>��o���y�r��}_컚�l8Gy����ë��2�������4g5	d���k�כ�@Y�K���v��o|�vw�#��^}z�iw�����z
ƞ�)/
 � �w��^��sot�Ƙ3���M5�� �O�("�p,�Z_&�ܠ�bOj,�w��.�*���\��S�)OIyx��Ý�Ƈ��.��`�n�*-���*B�P�z��;e�[ q��T+  pp�'H���s�p�@���߽��1
A�i��Z�$	ꮅ�=`�S��B��OEzM�w��r-�5V
�h��H=�Sd&�wzs�	�2�쩨�Lؾn�"+��xw��G�p���G݊�XXH��8�q	����An癠�ӕ�f�.��j*Á
��S�(f�A�q~��a��E8�]�7��[�9��ؐ�z� ��PP�UQ#@ӵ�F2���]�o�tH���cm��{��o�%{��"�;��^[HHPɶuK�)��ef�+��~��Qk��2�]c�p�f�]��y�_sE"��&r�:k�������� �<��ڜB��{��( Ղ�^��yP/�
*��K�����.�� IҎ�;TE=����CK����q�C��e�\�Kl(0!<���ev�,(���Q0cDȰ�7�������Ъ/�� �K�������;��s�l�!\�
�W���U���@��<yQ�nɡ��?	ziz��ӬE ��������[����:���j�(|����0,��_���>˶�t !��x��>����m�b!!ŉ��rFo��X��l�)���Ka��Rp5p�.r+Cn��g��?[g��n�'�<<���P�Ç�6js:P�a7��4�t0�� ;����@�X���Q�p����kv�;��;/��us+˶��<��sO��9��Pq��|}��������e��B
���zq �N�����5�D �n�;9ל �ĭiˇ�z
"|���w��3NZ�S�i����6ju:�n����� A���F�}KT�0�C@|�ڏ}큯����/}�����+�uL˴Lk�W5���e�c�dsö��ŉB]���i|D�@X����pb�`���{�*5P�)ks:m����^x,
@������r����hf�x(~��~�mx����q�?��io��cł��l�1o`��p{T�?0\s(�ʯ�SE�^\�E=  ,ہS9u(w�p�������D����Tϋ	ZO���P.x3z��q��[�-�x���s��s���}�����#��q�SEH9�ʥ�һ�k�L�հ��"pI8�i�`�Χ=	��$0��V�Ն�~}������Չ�"�r@�u��>�w�[o�r�Xr�w^���pkZ���q�SEH@�֏L��N�6�sq�,W]"bY=r,�M�ԝZ�<<<� 	|!o��=����E�����P�y��A[}�����	�D�QD��?����?��[����T����A5!��p�p����`<�fE�^-�@����8U�OOz��<<. P4�쀩[�������Oyk�.Q��7�7	Lp\Ǵͧ^zꅷ^x��g3V�Ꭷ�<<���H�K����hG�߲*6$�KK-�l.d�^;�}0~���K��A3?���� $�T���n[��t�B{/���ˋZ2I�tK��'��ﻧ�O�����mxw���UEB
 ����M>٪�O��Z
g@�\�7�;z���h!�ɫ�pB�I�&j��f���y�����F�kp:h:#π���O�~�
��O    ��xr�����r z"���*��) �\���ORJ��&��'��E|�w"�ͥ�b�{#���SǦ�m��!��"�］���9����7F��>�[���%g�N��0Y�� L�����6'������ʹ��L`<<<�$jR�P�K�G�����-bsh�"}����X���xǾ�#������W>�w�����iGV~d��׿������^z��n��頭F~VӌC�ڪHCW��=.DUQD(��x�NOY����b����w�����XBjR  �c�1|���F���;6"��L�Z 'f:�T�;�������,9���"P�����?b3�AX߹�����/�9��h���`?$*N��*N#���_PE�L������o�����IM�D   �a�r`�P��X�͓��T�hYӵ�=<<<�v#�  Aw�w�s�5�k��C�K����`1t��$��(�U��h*��)���XOrTw=�<Tƃ�s����oݶ�1�8�eI޲zK}]�p�R���!��ks:h腱}�g�L�i���1�񍾛ݎp�':��8"��"��.��k���T_�Lˮ�$���X�� ����+��r����6�׵E�⾌� B���&B�M�N�G&o�M�N�{g%    IDAT�Y�����E@�MJH���� ��^KL@ACP+�X��{|�"Bx$�V��Sh�ɧ������ĭ͍�ۡ��6�� N !2@��8�+1�)`&�rw�.�5����x>�M�yxx\�,^H �K�D9��b&�&޸!ѽ��l��|̗��L��ʴ�˅�I����)��d�7=8RHZ�Y.�����p�� �.W� +�t(��C�̿s�S���C���<;�8aD��׌ ��vF���E 0�����;彭S�dp DA�&9|�����S��'��Qr�@�$X�ϭ��������Y�xxx\�\�� "�\�dvb��=4hG����-�TEpF@�Z��3���=U�'����^*�'੨e� 8�ZA��Z��_փL�3��/�kd���+ƀ>������ɒ����8�>�����@OW��bS0x�V��t@2� U���ܧ6�*�;S ���v���uy|�>�2�����]��l��OY���q���R����蔋��d)#1ID��*aE�� ����1�e�r\�&��UQ��u9  )
�OB���p]
N���h����v��R/חy�?���?��ג[Z�{,����DmNAE�qU��3*@LR�nu>�5�Ɣ(⬮C�ת&n���ǭ�Ĭu�ܝ�=c����GD������tV�w�""�suG4��A��E�3  �E��� �+F�շ�X.8(qh���W�g�$�֯s�����JA1�sr.��b�5#���џ�X�5��{�������Z[��k�Ə��ck�/��F�}�g{� ��y]}vGwt�l�^��3c� ̫�qሂ(0���rc���^�����BH��|O�+�h,�%}��[!p�%UQ� �v�MO�˒��{�,!3N��Ts:�A�uu�M���D�29��-�aϜ*��Z�x��1��"a����u�Z���=�[s���ҽ_�y�͜{CR"6�DQ��c���I�k�>���m�q������U�i�Eke����;����XS@ �%�d*����.���R� (��=���(jw:��&�U	��?	@���h�I�*�BQ
��7~�L��]b[���.8K�]�tG8=vZS������E]싼�>t�[��^䅺T�2EVR�TY/]=m���f���M<EA��+OHy��CK����]�v����B
X�F���A��������?8�����r�8���O�8�7�)B(2�3!�D����Z�(�պ�r�,c����4%�|e	)�2������o�71V�q����N�����~�La%'e��ZgBU�X+i;� �L( �jv��"�>
g�S��Z|߬�jWs� ���9=w���3�:b��շ���ԲA�E>q�'��QEV,�Z�7	+��U7�2@ �)�J����?�Sp���Ń ;��W���y(�%�"�QP����L�#��uq��bX�+���a�x��z�E����H���mN�N����Ɉ"���Ŵ��Xٲ�J���7\N��9GI�����}A�dY�ӡ�Ž(����@��DĲe����r�t9_�;�$Qj
��|D,[�x9�,/�U c~In	��P�9^�'���\H(_%��g�Ҫ���7mw��D���wl�^y���'��DT$�1V(�{�t.���͚  r=A�e�a��ɅM�-j���d�<X�YMP$��� /@rA(@[��tp>Af �%�(0Q[�ޙ�D �I�����v�#�� @�I�����rc�%��V�D ��B���`6C��<�����nh�ڂvP)��c��T9z4y��pt2[4M��E��P�a��5�6H�A;�f���$��l�WǊ}�t����"�%���ݍ׷HA;���<U��F^9Q8:�-Fu�O  K��k�w6�A'��"�n+)=z$y��x|*S0k�������Z�ΠT
sM[J���ȫ�h����M�jT:CNX�1���d���t��B�d�`���+r �-�]�T�3"c�2"��Re���4OH-'�	 r��?<��y�b)4���G������ޘuĊ:�Z�va�f1B�(*Go��cA)(�)�bEǽ�n\ �8�`� �Kҏ� :�ӯ��S����-�6�K��|���;c,��1��*u
��l����wc B{,��mwvX��I�q�p-�w��[�~|L�U�HѴj-v���xg�����[	š�	w���~ҫ���hٲ��@��x�s��谚�Ss���h�����q�aݱ>f�#����;ڬ�PRf��.�9�����x⧽ʳG��jr�v�B��l��Uo%e� r  BN�m��5u����y|�p��B��h�-��-��"�	U�Ķ4K[��O�i�8:�;����:�� @DY��U}Y�D�-#g9��m��3�jy��ԥ�s������Z��eA ӵ�9�_��~���n(����]p��y�}B�9\�y���>���
��VNt^���k�Q\�̔G��ot�l�2Ӗ�]��k-�H�څ>�<d*eSM����T� '�D�Z7� ��]xp�@����j���P�KU>7cBD�/9׷���&[~v���m��W�k��+Q3��I�u�c>�����[8m+�)_��r_g1�K�ݪֱ��@RǾ�9�_R$�ڗ�k�dW>��	�24G Đ�egw�dP�7���#'w~33�Ơ��ZXU��J���c�Đd{w�DT��b�s�N���5�ZB���n�tW. �&g�
���-nDm4y��N�7Ow� `\�lo޹J���P%��b����=��	�����R�=�(������J� 9S:�X�G����݈�f ��x��5eC}|�*�= �$`I�N����F�d2c���V��خ���v*1��2.Ч�u�o�������A��;������X,1�mp-�gs��V�]���F$�X�O��Dl�N��Y	��B�Rqf�u��jp�򧷮��Z�k��P@YM��	�^O�ߕ�`�~(7��L�!PE�W��\+y�J��;�*  @���.���ı��`.5�+I���vkK)z�UT�RgZ�"���2�j8:�H�8���@�k[on4�J�����ti2 @&2s}<��u��#��dҝ'�,�w�o���Q��|V�� ����:��\w��xo2����J�I�mk��4�9?ӪJ��3�(	ƚ����6ND�O�x��`��!�����ƻ6�74�M�q��Ҳ� ��M��M��Ou��Ɏ�3_�¾����!k�M݉�w��$����"  Nx-�.
w����~�rs�= �y�� ���+~�:ߎ��N)� � 6��� ���⡱L�<o�� h2[�(vDJ�����>�A�f�r�ǥ�l�c4�6�H7�ܑ��S��	rt���c�Kc�$n!2�a���d)�zU�
�"L�1�ǝ�kLp;TK����{:�&�$C��P�39*����kMq3͝�����pۺ������.aB�ݹJm	L1t8'&�fZ�q�蚓��9��ol���P�/�d��\w:bT�n�Кi�'bӭj\3ɭ4�s�*���2��<���9�FP'�;���P�
� E�g�:�U��oLLܶ�7�+d�	��qo���/ ��c%E*�T]3ͭw�D\�uu��"��|Ξ[�DUeO��H�9��fJc
wʮ1Ν"���������p:��1���B��Om�]�d�B��L&���-�Bqg�d]0�E~v��L��ex���eADS�����bw4)	���"��#��r�+Ĺ�}���B���c���=Z۬lHL*���D U�p��:&�	7~����ё9G�	�ahB�s��
C�{�^A��՟.|��o�g$��J �;|Mw1i���d�Nh�� �RZ��7f�M��Y-z�@�bH��5��)5q4+�W��_���?�&)dQ�Ǻ"y�9D�Đ�x���-��IA�<\�W��[0�Z������[�vH���uG��������@ۧ��� E��_�x�8��[�2Êqm}�ӂP�Λ�"��*R�*H�&&}�w�����c��)�G�O��Շ��u��w�3{�<���a�[�V{H�L�����Oi�{��]<���X�g{�[!�x��⳷��y^�vY�VkXrP
�>�k�W�_ˤ�S.�<S��S�BJqk"�K���:V��H�+\ Pk�=��|�p�8�O�R�g��!���=#��
���B7��gUA�����]�Ĉ��Rx����j|��6q�d����K���Vju(Y ��w��l��sl��R�/Y�}]�c��U�	�9 g��~�;B�_ӕ�?�f%"!H9hyN��ׯn��ձQQ��1E93�/	�ֆ)�D�h{c`h-��TY*wN�K
�_:�&k���؛��; �5��� ��'D���\��N}�����M���*�^���Aęt<Y�oE_2	 4%�D6J�չ���sɝ�I@�
bcD)I ���@�á����d �z9�J�l��}�̾%2�I�Ê/c�a@�����&c��χW?.�*��F%�Y����7+���<�YAE�2��C�����	�H���Ъ���3�j�B���܉�n�~��	3
�4,����� IwQ:��~Lu#VZլD�H�չ��nf�A����
�\�$�n����`����/ʑM�D �z)�Nm���#�:C����(P�Ϗ%	�-���$��;����\L QkR�;$g�����o���U�׫_W��EN2 ��c �#�g��~�aJS�����I�nd  5�+�r�o�����ԯbj��Ny�y�R�]�U���LA��H��.mUlR`��������ux[4NHӟW3~���`g��S�|k�"��`� Y07%ҏnn�
�
�KX�l�S�j��O�%��m�í��=��햂kPP ��)#��>��>�2�Y@�v�cS�g{�#�y�e<�Q�#[B����yHL����f2{������ UAPD�1Y�]Y�u)�L�p9�o��S:e{��UD[b" �k�
c ��A���Ъ�ʁUePi�"��{\c<�3�U�$AD`t^(�LDE4� �ѝ�5�F
tUT��R��t�]����J#�<�Ѕ@��D�d9�>��y98��fB��w9��]�'+ŀ8Wz�@�� @�)�=���8g��Z�mvi��༤�"�8w��q�r���`��R���c%�|�w:椕?"8�Ɩɖ��c⊻?8���,���#�Gi1�"�9}�*�.q�.��]_uUԚ��< &�}�w0�Gd��-��M�u��z��3�,���,!`�7v��'J"��/7�J���-\)_��X�j��C&��"/0�2�^���P�A�뻣[fBae��L��P��O U2�7dnY�x���??Y�ܦ��L����+">V���` .���;A� nX��v��x�rxS���v��.��N��(8\:�?;�30a{�Q�EM��-���y�ǘ�7�Syʱ, 9�A5�]t�VQӡ��V��4��c�����6��L
����:�s�L
i+���1�B�<^��Vb�����5+��jݍ���l+v" ��T��(�Mx��#Z�-�����ת�"�R@��A����*rDM\/w9����!��Ā�pۙ���CŴ�-��Sv�I6�7������!E�/4� q�-R�2�~o��3���W�`�_�_h���dcl]L���RK�'�.K�k�/5=�6������ע �m)O��B6>}�m �w6�u���l ���=�t��#jaws쥣b�XXH�����������|��w��4��H��;�e�@����J��?:A������. d�9C5�Ԅ Ek�c�+���PD_�# X�-��O�w�y*j�URX�����¡4��v���n�Z'H�JX�@D(����yZ����j�P���*;�n2A�396f�`TiUx��g�C��9�K�Ho��X�d'p��g�ڸޖ������9UT&���[�cϻcO���M�п�K��R�#�Xk��Q3�icD���E�l�� `O��F��| 	]I��OTT  &��f�-V�� �)Q-q��(��������ԫ��T|R�ώ�|�%���΄��U�n}- �N����k�Lx�RW86w���o�Ml��m��3��2t���	��lbi�wh*���+��鲾��+N����]�i�^ek�Qw��LDlL���Pg�i�ڋ�9-��Ҫ��x"��\{��D�khմ�Z��*.`��H �E9�	u��R����Ϩ���QL%����{B��1�h���3� L�CׄV}��|/��T ��n�]���r'��. ���B�@�p�hY.��)¨*&CND�(�6����=��2ȵ\c�4������b��@a�V��;��B&V����o��B(( @��Z������pʧ���z\� �ulbj�T8����e��bP5E H@�ͦJ����I���|2]���g=. rM��O�9�ぜ�i�J�2�� ��t��A8w� ��I�LUy�ഴ�n�����hq��Y�����e�48w(�>용3_a��!wKf�(q��w�I�LN[p- ���[�>rM�},9NyĵR3C������=D�^�ώ��7���F M�TB�`7�*JE�w 0��O�d&U�&�'�.OPBQ@����w?�o{@�cn!(L
��#S2=��	�0}�Ӳ^ց�Q0(3Ab"�c��/;?/(��&� �D�Q���� �9J󧸓�ku�V��Q&Gf��JT\�82)w�;Nypi���G �E�x�~���ڀ��k�E��XD$�����I�T~j�\0�F]$�����̝j�M�LZ�V�8��.�UhA "Fv�H�ie+�m�dq;�O���C�:V�M�!� � HvN�|�HݯƯ=G q�T��S�%"�q�⾈D��S0�o���Jt˹�ܲ>�����<(���!�v�<�+���J��st'w
��v��N��0N%s���1���9��w ;K ��ד�vJ�`z����B Qrrr��/�����M�ʵ2��KV�#�E��x�����T�9�G�l��Υ>�<9c��U_�m��{f��3�19����~�h���;\��<���q ��to��Sg���m�ɑ�����?{�gWu�}���9��ަwu!��@���bن'~��&q����8���q���M��1Il�6q����&M�k�G����v����㎄4��Ќ�:ߏ>�H���Ϻ���k�������B���j�6�>AE�J	�����/�L��v�C ��1Mg�H�������G� ���(��6u�CDN�3�� J^5z!J* #as3U��}��a�N��>A�;\�~�`�vg�Y�)5v	�>FĹ�*�<^��� Is�w���H����J�)u�� ��
&y��V���H��1��d�{La���k���~����{��5�����L�0".�|��w��s�h@ X8^xG�1 @$���\��(��L� �#�R��o�}O/"� 0���&1(H �D�.�w���ǽU��+�z��w��$ �;��8�>�	H��x�c:�p��a�T5vɱcE�*t=T���BѽXN��C�rh.9V�C�]2�SJp�.u	N�f��^��R�H���r��'��G�������HF��0���j6Iqj��U_a���9�Q�(y�+���*ɧ�.*�?�
�w��at��:���	�p9�����v鈿�}��E(�B��ܤ����~1Y5ݱ�2���)��ym�yn�|5W{��$O����ĺR����"p��]O��a�1�mw�hi#�WL������㫻��%�.1R���5�d l!����i�;��8=�|�E��6�<�Ҿ����rTB�6`$7��� ���I���ԃHc¸�3/    IDAT����ӂ���MZi�I[���_DT�R��ڢ����� ĉ�k^�4�J%8bcA��eK�4�c�|5W{"˙p�!3�����2ĉ�d��J �BI��z�:�٥�'�����%���u�m��ˎ�[�"���܆o�.	L� 0��m���C6�����13;�!<=f������
�
�L��ML�	/'D`��$5v�xKd�9� X�I�*�Z-F�?�P%������.�\�t6 �sfj��k�KADI��q&SQ  `s�+�>�YR�U�!'o$_�2[Q��$r��k�H$���4��� �`s�3�ڗZR��ze����Zo�v�� \'^"� �����4}ܞ��;3Ç2KC�Wv�ɛoY%�0�)	^Dd�H1��ny�p^���u�+l�5�׶�xe�켙�`�v39X�v"^"n ������TF:J�m��	6(l�5��iM��Iv�H�4]uP��ӽ�Ŋ]�]\�Kqww(��^ܝ�R����Cqw���7�˿�'yv�={Nf3�5md���+%�$ S��06띣x
��>PhtѕQ$W^�di�m��$�����H�����tS��$蛠|�/���Eb�e�Y�;̬3�hA:s	��n�H$N7:��R9�Ϸ������$�7ĺ�Q$�>K'�� (^Cf\�P DFBT��O�_Rဉ 	h�/C^�#�9��.
�D��䨜 "�?A`��頬�U��o�  �Q��9�A�ad��_�*� Nt���L��H�Y\D�ێ�� k+�)�#��QE<j�HGh<C�xJ�u�����Gc�($  ���q�~1,���
�^Ľ�p��l��!��<�c�ugRj��Od�7|�(��Qc��$���w��>��4 p�Y:9���R�O@�ؖ�)�� b *~ �v�������uYݏSyth�ǣ��O�=9pצ�ޜ<�%T9�������ý�1�Fz����QF;%��w\���m����ƙ�k�����%С�f�������#�GJ����P��A��ӛ��ۤ����uWW�#�4��u��+�M��l��;��?�-gO|�������|GG�P��G�ڟ  QV�T=���P�q��G��P�����[�2w5L�zd�T?̌E 2��`����T��G�VΌ俹5!k<
w	6�}�>��=z��K �v�R;�c��i�#�cW�S�;����`�.p�Hŝ����Rϭ��Q�����E\;}?Yݴ���"�!D`�
��WM��޺R����G2=\�FI5
�=l�=�(4�X���`�^WE�v�#�%�A����x���J�qel�=����ռ6�,X#(/5U�L�� ���n���9P8)j�u;Ð
H�����8N��I����Q����4�T�Mu�~�M�6�R T �	O�O���vC�c������ѺF��*D!��i�`6��~�vn��KS���M 
�����x�_�|V�6�#�~)�U�EᘞOܜ��h0b�uC�� �
�>�\k��X�t8��d���x.��7�OD�$ �B�'���_ҟC�8D1��y:���ڦ�q�gݍy���KH��9�_�zz6��3��+��7z�>4�0�>����hIX�,/`{;W5���Mvq��@X���){lL�Vm�;���{�����@܉Ǉ��>:!@l�Ζ�Q��bp�!�A���O����	�t4�}Rf�X׺��������֬�ۨD���`p"��s{��g�=K���P*XK������}���v����9��� ���m~J��/����/��H�5�r���8�G#w�w��ϧ�vl\��Q��I���$T�$��پGS���"*�Ԑ"���/m��OzZ�M��8[#3.�bm>[!����;]ȷ��ZQG�����a��� �Ь޵5��ųS<���,����m����_�ŉO�����`Y���M/��s��J����M��7f��ߍ���mS����6�~�v2b�q(�5>n5VB�!�3���C���Ϋ��ߑ�����K����[]�X;�,Ο��Ϙ�(�qg��`C_����k,�<�����i�?2P5h���>wX���xw���&G |%]�wd.�	�A2�nii�����ʯ�RU.�BM'�ˬ\q ���[��Ai�gu�x�<WX�~23xx4?`�9s5����8��w8q��?XyNlc���?s]�"$��`�#���?��}��_p7���1Ɉ��U�z>B|[D�HhW�>?���葱'���u,���jM]��~$25E�?d��j #����U��p��J9؉!��󇥔eg=�;R��8�>ʲe�m�̶\=�m{�SWZ;8ĳZț�'6ݺ���j�\�u���g�C+�Ӌ�)�B��0�Zlk�~�߿���XҐ�[��w�C�P�����J�@�v�0��cxR��Z��篔�t��Yw�8��Lv��h5R������X�rc#�:�<� !cj�*�w���p;�_�b?;�4ͦ�mG6h��-��˝V���)����,��5����>����mlL��D�
��H�	1�:.�-�0t�H���/�C	��jN���� K����t�F��f-B��kQ���q[� �xzϟ$�u���ԴsRC ds	R����c�QjD+�/��8��i�կ9�.�/Bט~?~��fG�2�.�X�k��^�
�CJK%x�s$p87O+؂3��ܳ�L�}���Ke>��T	Υ9)�/�m�k�z�~J\������0q��{�%�����hg��yr�<���	�NyZ"�`�k9�94g��5(Y�d�X
B��!����[�(���S���e� �<����s4r���ɡ�;6�"ɲ��Ҹ���MF���t6��=��rDpȇ���h��VN���o� 5O��~h�i�g�c���3�3���&a�/�Ī���\%��!l��'��GOWÕ �� 4�"8!��D�;`M\<R�QAjXX�쩁�����y���c�q������;xn���A�r��~��Qq�A�/�E1톅�Y�@�8-��D����c�5B	d�Ʉ����V:�l۴B[W��C���.Bp�3E�^����a�Rd ր������1]%�=Jr�l�ӚҤ��즅� @Yj�pv�L��ȗ�d��|�y����ˤ@9>���G&L٤1UJ� c�|�$�~�_�;r�X���(�:c�d{������|ȉW������E��X@��> ��i`�Z�w�n�=H�J����f@@�����Zg�h���02��9�X*$=q�` g��o�;�C�o�I�n 8�k���HLV:,P���}��kw6���z��Z<��'��5��d,x@�IDۯ��}YG�1��l�1/�% `X�Q2>δ3P@$@�mg��=���aH���e/)�"6s�O�/��EP����q��n4f�H����6]�.w�w�~�p1��y��x��֕��V�t{���6�kN��r�o|�]�9��hU��d�Z^�\�l��9j<�,u00P�&��!�/�!5>Z���y���4l���в�� ,�yyq��S��J0bö*N߬�O?�g� ����TD�aoJv ������'��y���*i�أ�Ƨ�ͯؗod��G��a�I\P�IG/�e�n*]���ئ�qAb�1xl�I�~֎Z�j�<��e<4b|L>�Ch�دh���$N��U�-isM-��>�w����0fG�À
8�r�����-f�.bdU���H��h9�"�v�ł6��˭��.#^J��>Ji7�k3#;�z��+aĨWy����;��3ݓ��dεkrHb���X�0v~���k�C�56��:�������Xc��yWn^g��c7�������F��Z���S���;_����X���D#'U��M�j�>��?����:g����McI��i8#�y��Op3������ܜA�hDt�U���:�@q��
/f�zRXg�t�)�GE�H�����SZ�U>��%��-=�P$sܳ�į�3�4�z9k���~�Ɋ_��65@c��B�f(��56�%���V���y�:������1�/�� N0��/��e�M�_@�u�n��U����8�-h��=��G)\S���<`����\�H|�����V�M����U�RBv+%Q�{L`��$w�L�rt�$uV�����|`��x�;���u��~�y�q
V1	��x��������o�W���(�ܢX�T���lJ��)3ʩ"��[Dnڜ,obwY�LD��F�Ąȕ	h�W�+�=S��E������K����b��
Xm�S,�X������v�~
%�k%��œ�S����(
E��4������s�%~���m�_���}zY���p��s=�`����a���K�hmT�����A$`��E��%�WhPR���׷g�.�i�(��O�ROc�Q��� D$�݅����͖���� \LY�7Tv�_�\�2�4��=j���E
m���%a��7 у$���?8GT�F����*cK��*��2�]��SJ��j��F�� pd��k�JN�Ќ��|D�?|��2"?�[�%
�ŝ=Ef�k�C � ?9�@H�r�̪E�,8�e�!	�P���Gѧ�X�J8�,�a�/�6�Q�JH,2}��AV����R[���0G��1�P+T�����s����#�� �b9����T�1�*����O8�S5��|�8�D�c��w�����m,��!�Δ?m�r�Ur�eў�Ց�6>����-ŧ�?Ѥ�[�C�\ɢ�&����y��mO�6gl�W~��Ei}d�XP������T����=�	d�iZ$[�:�7e( ��W���ߤ2�ұ�l	N�(AgNJ����o[`@����N"����l�#���&�S��!C�a)nfH�v}���j�'DA�D�歺���`��<��k�:JZ�	��QF�nz��{��acڂ�o��Gbl�T���Į��b�ޤDhqd��e���I�sJ��U7�fN c��uDA,��şs�*��p��KGO�����5F��(-VL
��M*��'�/�t�pjs��T�K�;��ÿ�)���vX?��1�i�L���C.2��h������
�?�w�)��i���a���p���wey��)UU���.1݉ɘ/����d#�m<��2�SNo�u����������0�ڝ8^����gd��{_�f�"7z���6�O�]A�?Y��H� �}�oD�o(�I��)��8��MS8�S�H#�2�bt*p�+���\���"�26M�H7��g���i�H�}��fz�ϯ�Ў��w����g��|Ak�qCqF�Y�z;Sβ��Y�I�0iQ��9�8xZ�7�B"b�8�ٝ�%L^A��S��h	i��VF��C'���D|�I�O3p~ݱ�P=i���C��"sv�ɘ��"���ҧ�0(��T��	D������N�*��c�Qa�YF��s�;�؍��Q��Vud�H�����D� �����RO�Hf҈�������ar���>�p���
����p�e��Pf���`����ys�j�	}d�t-���>�'9��9�+�b�P�q_4�7��x��O���7�����R2��%t^1���TL"�`�����$�L�q�I�{�)��W�2�w2�~��۪cj;,��T[H@/���������ICC�pį��.����i?&FB71�XƮ�U�U��Z�L-���EȊk��{Kr�}M��4�#INh�F�+_W�$!��ud���寉;��R��d89�5�q!��R�Zy�ڣ�Q$�k1a����ҳ	�b��o
����T����9��������OS��}���-��A)�AŐ���M8]@c�;;�^l2�'Y4�N�SC���O$�kE�[��Hf�:�e#�j˖�޿=�V!K�Ԃ�d�~{�Ǫ�u��s�7��.9ь�00*��ӡ�������~�D9H�r��������p�R����.ǑQ�>q�U�214�����6,V�m.��z�R�R�_�$���JKM��՞n��6��zPmV{��q�_��kHU"R��"EbMh���;���on.��T���w���&�S0�*33��>�H��UU�X�גP�C���mC"��K���EUq���G42��M��n4�'���/�c�*������39�L\�Yʖ� ���
�a@c!��~&���^b�@P���ةͬ�P�g��<�C�m��5���ˤE�Sֈ�,	�q��pѳ~=��:^i�Kr�'ߊo�+[ե���o�^�Z��<Ti�~�G2�� (8�&��B^Uz�6��QQ�B�_;U���' �}�C��l�	�c�n3z�'�8��CZ�M3�8�R�}]��8r��ؙ��jg��|?�^\o\�+���b�K O 	ʟ�tw��%!����|kurEY�b��C�{�Y����5�k�#����-��G��חY�g)��:�#������	` .s��%��7���Z� R��_����-/�:���mdL�󇥺Q��ZoZ���SX�W�k�ԼÎ�����K3�l�\��N�T��,���!)��0p�zߵz`����Mm�_�����]e�]�z���3����=��&]���§엍CW׳(�5����l�2�N�8��ӘF�1�zM�W��~�loa� T0�A�Ǽ�i���_�ݿ��ѿ_Ϟ�c��\�k�J�Vw�'Gܜ����~J�l�9?�;�M������WD���Ql'������T!aPS7� ֣R�p����FWDf�i�aB����U_%c�Mf�\��V��Ku�����`i@>Jjr����h�c���I����0y�V�k:˲/Qb����s��u|�ݺ7sO�����[��Q�r��n?��L���ǥ6Yj�,:�v�Յ�j�F`I�Q�#N�Tw��Tr��=�_�������n����kr���@���s�"�jBf�m`����k���ո�|��3/��8���\�ӈ3��С)��d��0�cB
��c�\.��%�,��7�^��!Ė��,]�^}'��O��(
_��~�V�2�!@4�2�3�,��%��	E�Mb��_�n�t=ϖٳUyF6}k��|_�m�GuR$�yM�n��Z��������.pϕ�� b��;[0Z}���ϒ�,��@gR�VJ�d�,!�����v�������k��ጀ��n֯��Kk����u���IG���=f�KmIRy1���?ƿ�.���HxR<oMI)2��<�C�������Vo=A{?��kɲ�4��u��� ��J�*��I�\�tJ'�^������;;_\ W����_�̚���QIy"^��zw)z�y���ղ�/�)l��1��E�����lT/c���h*e���UҨ�X�f����15r������?��Ƶ��U��X�q�7���G�-�Z�*Ò����/������GԱ-_f���t��^�;�0�Q�W�x��ٞE�挆�J�&?w�7(á��w=��%_*��&KPvz|�����28����Q5�T4����u�wJ"7=RiG`=Ql׺
�2�����\;��BN=|tP�9�Z�գ�G+u��þ8B3��j?M1�k��8�uI90u���؉|$�1�T����+�)�,����jJ@���p�=���(b��UF�b�5s�H.�2�P&�	�����ӎ��6NƏn ��sಐ��s��9"��8v�NE��Λgn�幢�+e�p���«Jr���R�8̮�������� �(�ƻ��ws�![�^?qXUIm�>D�L�םs �-����]��>|	���}(�s i{�3IK���kwʮ�� ��ôB<.�0�BTѶ�`�C{|$:�"�
J�����[���$��>�J�?��Ѫ�+�5w5�W�̃wÏ��C�䏩y���G)�6�}�z����$S��N"�6�HO��5k.�qc��-���$a�w_e��=�H텐ȡ'��G���"��%!ֿ,~*�����q����ܬ${�^r4a '݇���r#�t�_֞׼�R�H�2�q�9ݿ5-��\0��VGݺ��O[���Z�TDKa���k��P��u���~^����ǆq[�~>��ڵ<'�ߡ�Leo��/�.l�< >�N��}z�:�=�T�Ѹ������[��n��՝�:_������1^�wA�L?��r<]w��U��k1�(8�N��+�3�q�Aֳ�[���k�����w��S"KdKڧ���+=S�|�͟W��0�á�n�tґ�IǗA"ܼ�Z۩pkv;�n@n֐c���$6�Ǳ�CB�.C��2o׸f#�^qJ�`�������*������fҹ��U�B������e��"��SJ�Q #���ǼMT�o���f2��6�� ��+�<=���B�w3�z��|sp�P��C��a�Y�{��0_�YѪ��9KtD�s1��^|N4���[I��O�(�����/B/q�Z���S|�f7x�,��p�����d�ܖ��f� �6.W�3��~�������b	�iJ�I��DĦ��(#�2�%%'��]a��ԍ�L���i�kHNך���&Pڀ��ҕ�{�6 ġ��6ە#�`�B �0���D���(`������u�E#+4i�j�V����K��61� ]��I��u��A�7�*	bOx>�A�����9`]�SB� �l[N�����?�O+a�gu�ݰ��^��>�ވ�������VyIx��c�&\���ؿ%�6�]"�f�����'���ҋK� �p��e6�I����]6�3��梄�ώ��a�a��4μ�$��R$7��1�Ǒ���c��p~�p��Es�P�����Z �X��m>uB�V�|K?�b�Y��ёD��QiWW|�=�bx	��ŦF���zj	�ˋ�uKa�g%:m1��S$:�����W$�S��w�W6�0lC.Ur(��|`N�ú��4}�%t�rk�A�����|�ҹV�����k����&����j���Cj\q���[��{B��L���ì'��Ƌﻵ�K�m��x@����E��/�����F	�`�����!�u,�w���LV"���*L�8��A[65�%��o�z�&����  �#9���S�5B q����w �ݼ�WX?|[DK�@J[QѡS�;��.��SY�O�@~[�o�+��-6��!&֫]6ct]?��S�0�����"q~Z�
��I�v��7-5T"È����VhEYF>֨i����ne7h�P}N���"���P�U��O$ ��h]L�g��b?P<#��iH�bQΛsDz�&]��l&J�������uT���y��d���u�J��~Ǽ�oo��4�+� �??Bϧ���F+�,@��C�z��/?["��`hY�N�uLw���}4�O��/B�����Z�݈`�����=��Bjc/_�d�ń��Vy~��nk�눅3���β����e����3�>]�"�|�Z�����Y�&S����T�Qv�=�t*sG����,2$ ��Hyj˞����^�e���K�z@7�vN��xG���N�Fy�!� ��ei0�����������(#�8y���Yx/�s3�����@����LP�d��hv�
_�),m��A���~;T�&&�Z��)z����0��4�n��Q6	NH�A���n����!Љ�e2�!(�F$ޱc$�`B!�W­�U֕�ɉ�>Mp�j����Ҳ��{K����a�eV'�yG壘ty������ ��֚dl�P�z�f�m2�.�i�@nֺ�gT�z�cI?��CI�E�agvmy�1��b£R��<<�<��ʭ7��1636g։M��9z��0I���6<6�._�<����^|_V�O�
��=�>Q8bwC`�\�G��+$�Ϻ��S�<� ԡ��6�8���7��j��X#��)��$�/��*�iѡ���.���_��, i�h^��tr�5+��e��Sr��G��@t�+J���.|�Ahob��`�� ���~ƍ�����ޛ�-	P�n����LL��帵�\D�H��`�\���_����A�N�o��o�KJ�{�^J=�`��!���4�]��]"�9[9�67���W�v||{�s[v�gmzqF������b�r,\g
�X�4�n>>�ި1}gW���l�	�ūs�q�T�i����ɋ9����N����Y鍐���J�Ol4li�0E�R9��O�@'3��������&�^����G8�%�"* ��M&��"{���63��X���/	R�K2�Z�^��-��La���lڡO1�!�8B)a��ŕJwR"� �P��4�V�D ��3"w��v�`�v�}�P���w�/.��=|У���Sx�%F��9��NhGZL�>}w�B�g��k�pH�Q�j�E0W4&RqV��� �pgI2�o��ճ�'i�pƒяI�]_$�P �m#���ZS�e��]�y��C���Wl"�i���H�ឌjq����H�% B��o$����`xu�ʇeH�cRɩM�qJ������hB�A�'�m�T��0��mA����2���⟉���@c'OzU�8�0���Ç����Q���\H���z�W��S��块��V�UF�]E"~��x3����!��z���S��`�*�lu-Ͼ�w�-Z<{)�%AR����K�I�M�+���;����:��f�~�A�O2��	�<�Z%���~mƿ9�P2�춮<q-7.ys/��:)jc!��\@Վ�.�m|�dbQ���H&u�$��}J\t^R��f����7�����Ȝ�t���R?w�$$�*Z:E�4/��B�𸫪��98N2�GQ���S���}X;�9�ۋ,��QH���-�T��10�̹/����֙��H�%Q ���ޜSh �r�e�i�s%�h��G '��L"(���5��v�a5�N�[s5��X![%�[��	2q��U���I�����֒�vxH������$"/r���h]�B��d�W�zִcȨ⅐� 	c�G��f� �,���)�C�`ɔ�x\-֫G�I�ǡ�$p��)���A�K�s�j��s���%�	�|���}r�So�p����:N�� f`��[��)K�y_h�ҕ�h=�9M����:�f�����Æ�bE��񿞣�r��\:�tD<�=9J�D���m��쵷��4\��A5����Srf4�+��>P�v�=gj�Wub���[�����rb�6���?�&���9My�3+H�S6�����g���X�x�}G[{�O*����Ֆ���v4x~�ӟaT���pb /We���.7w���c"����d��w&,�w�o�w_lll��
�Fە&�3OHէ~������K|c�
�1�F{����'��f-�z�;�Z�-=��}�T�y$�l+o��Pw���� �UI�!����#_���J4��
{ծט<t��Z�I,"�Ǡ`�ܘg��F�m%U}O�hrȕ�QyA�;О[�&�p��m3ə�J>Mqt(񂓀�CO�#�(���� �/��J�}��!��.��#�6��
�(ˋ��k� OFҶ��^�)T��tܞ���001�V�;�Jn������['��@��+��G��S���s��1�vbQ<{��x`�<x�mmV*c*1K�l?��j�iҕ����@8�4�h{��v6�.���&� ��$Ft��w���k�_O�xO0Ǫ��vB�;p� �`�(��.k0�x�����Z�[M�R(�FxñML��_��l9c�$%h7�FfG��H(w��x��s��+8ҧoНG�ב�G�L~׌=Lդ���@$��_�B R0�Kq0��ʀ��K�,�xiF�n��)��f	u�'��AJ@?�����Y��?�}�=��p  �u$����5��A_ǫ�660�{��v��m��p�ª-�5B��蚷iq��-���u�-��Մ_TC���jq�P�!�m��bH�<����D�nh�sΌ��_ &+����
�T*e ��� �&7�۔�pb��jT��1D�Z��=NԷ�p�u�l6F%3Y�:[@�l����)��0u3��'�8 G�DZ2�eFH��xRا��CI4 �tOtAT���^�,��&g��\΃:���ڦ�=k[1>yO#O+򺞏�ٛ��m�d�5S�<&*R�܎Y��nƊ|4�#�V'  K���GQS���ܠ0��C��Ι���ǔ����Ǔ�0����(r�d�+�}� �����_ ���_/};�m$[Ұ!���/^/<�������`{?��6��Av������ޠ���}�b�W"r�஢ ���>$x=/ɪ{K���*)N���Ԑ�啖?���\,d�XK��v��3�m�˞(T�)��X/�Pl��0���5]q9ض<'�'�G��w�)�B���ٳ.d��nUe�ԓ�����7�Gݽ��~RK�_�'��FZ���V��E^I����6��0�t�|6��̅G`����ʐ�dzM�4�	��/�U����%��_�����+~�]���s?X}�,s#_�t?#��{^/S�kzn��:�W6�!һR�h>�'z�_�)ʇxr+"�v��Z*!t����s�ͳ72Fc����Q��Y@��y���:(1HI��$b���
�P��" Ҩ�VGўo��ߌ��Z��qr(1�}:c9�Z�6Vm����&�B"��=�j�
��"��[Q���ȅ9��'�~cL��j���M羽l��qc�pm��ɟ�ʿ*$:�e@��������Z��o||rf�yxL�;�S�Y7�\����O�徛*C܇sC��m���E��1��rmMe�v?��}ȟ`�e���q�3z6ܖ_��W2�i"j�=��:�j���Z?.��Uҗ�W�J�혀B�nծq�v��3�$��.kOZUi��0��"����iK$�,m�+OF(�</vv� �$ʿ��K�����9��u��q=������.���^��Z������'I�*F� ]���]�ω��so��̻�l /Y���l/|��񒭯�-$'�a����Zf�Xr��ܢ�A�Xcj���D#Z��Qa��~�ζ�����&�G��z�m�_��[e^���ڜ]j��T}/�M���
�����(�͋�$��p*�-t#%9r���� �7�p�T6�m���JB.DVD��S@��\O�ڗ�N�9�Qr1��i�դ��oI�ؚo
�p�s��~z��:@#�%p'�T�oMƤP����(Q�D�oFg��Tg��4�?�h�h�mj�m��e_��טtz��` �qxҞ�嫾�;"�YS����Ph��A�$L".i�"R�^+��Ĵ��s�]�k���M��(E�+U�������}rJ�o:w����87�u6m9�Y���@{�&C���Y�d��/?Z��EU�gY������~����j�R1ϵa��EF�#��dSU�M�_�)c>�80"�\��j�g+@{��Û債�ç�Q�*�dsCjE辗$~�z�_��-$����9�A N�����$��B��MĘ��'b�%j��X��Ё��V��������F�� @&�aj�uV��aU���Oʟ�]~�C����I�:�&��ؕ�j�B4��+�����,���>_h�V��H�h�)���8�ȅ���ͨ������t�w��/�0b0Z&%�t�=C2�hƭ���n�0��)����a�I��^��ة��Q����W���5}��7%�p|>70`r`0�^�xy��z6���������|���՝C:}u��|o��{`��5~���ƨU�_�GVB��v�9�)�o�gͫyh��J ?4��!Һ����`A�*�J�g����¼_�0@�_EG�����m|�W?���0F��6���É��J���%L(S����u��w��دG/�'q�z�C'kI�uW����ܛ�zUq�yڞ�z/e�z�7z��DuR?�h�Y_�Ja��1� ��-�B��_�Sk���#�J=#�cO�88�P|Ғ(�fS�2��m�?P�I� T b� Auҷ����&s�_ݒ�����gj����������k�ݮ`�1�mUo�Q,��bH]�~ߗ�C���Р��a��}U�����/���ﱂȇ���@�W���6�ߟih>�5��*�'�	%1���Ú�9^���5��w�9�{p��0����"�9 Nt��dF-���F�g{��"���Y����r壯�m;)E�����}?���v���-JVf���ЄBk��`��y����b'S���Gp�O���,@�������+�ex����yc�pNR�(�0b=��*++��J���5e�[�{�
 �3��]��a��z�D�|Zk"#�T����ؽ�n���6��6�ؿ_,S5 �;��SE_X�W��I_H{�G�H�2�	�-�e} ���崍:�ݗ�+i�8�\��<L6�K�n������m��}�'��8V��ť� "�W� ��A ��c&5)_s�=���l�����x.}���W���֐ c
�n�P��ť96c��[�#�;b" ��*��I�� !9l��]ͮ����&B���n��V!���n����v�z��lOEp��~�����8��3LC�'�Ic�n����V�Vv��zW�(�2سW��%�%�)�,"!�vN?��O<B����A�P����Nt'�:���|f�R�b�}��\r�̡���;f�<�6x^}�5��+8[:�;}mN���Ddr�hE&�$GpT` ���E�ci�	��Σ\�|�[5Uҥdm�2��>�{{�����ۏ�4n��-����r}��F5*w��ҙd��]��z�$vQ��R��ǉ><[UB~��M��%e�
���!�!j\T�( @t�h�+�^?�(��s�a��詟x���9�c�o5�M�N�imv����@��«d��<��E�7)���i�n*��_ZU6�A<3�ٍ�$�x�Jx�|���4�������,*����Ѣ.����DL;�>}�����k���R���y�ߌ/[�</��Η�غ�>���;��=�9k��E+p�X����<2C�P�[�#3A**����VU�GF N���sEa����lnY�v���wa_�)= (�l��8 �{M:�Z{Ni�9O�k�z�g�qG��}�����6m�H�׀D���F��y>�}�:����3��Q�=�<�����2�����k��J!���,mǿ�>XɎ�J�Yt��BX�k>�k�hë��#Sϻȭ���f��*M���C���Mч��$7_)���g�l��eR�� ��ViRQ��~��X��~�4��u���ؖ��惩��p�%ut+s����oG<�q������4��dv�6�ux��P���4��.A, �����<.%j��oj�؁#4�8N)����C[����||�
�̴�"��V��j	���y�b}��[��Y]���Cit_�|ȥ��.�վh�:�ʈ3��IZ�C&nr��yI�������	�[QO%�52��Y\�=��>-N���ivg��<Zd	�ahW�uFK���>����OkL@u���l�R�L]08њ��M�'���
 
0�}��N ����>r���`cv��E����M%+	�Dϵ��P�C  ��������n���BY��7��O>�/󹉃dJK�.]�_a�o�v�0�IP����Lp���Yѓ�"dv�e�z�%"qa��4�x�N�/a~���)�|���nf�G�n#�Γ8;^� �T��AB{"��e{�P��	~�(���	
U$�D �i�T�ѩ	2Y~�i�����8[QK�2�'����n�T2�)/沤����%!pr��Jad��(oC���,�$� ����3���¥!������2
sZ�G�-��jw��::���z>�ʏRB*�ԧI/QTt��&z��.�*���O�p qu�CA繵��X����.Q���.��W̸"� �h(Q	#~�\po�,�g;\�Ҟ�_- �x#��
h�Q%��*-�Q#N�Np��{C�FYK��;Rͧ�a"$\B�;��4��V�T���X#] �8�0 ��/ ��du&�:��j�z�|���QF�B�͠E�:���Y}�oC0x���X)#*t�y��ns?q�ҳ����!Rh$�ﴚ���r�^��O��F� �e[$�?m�9��8Ff/�!�?G�q,��T�:'�h}U�}i�S���Y*<y��jo1b��*��ߧ�d%Ɔ����A���wOYOƼ�.�>K�ƾ��?��q�~��;2������~�mtA���ӎ�����9�P�����sSOW��n��?�B����.?�jr��O2�`'�iUL����Ʌs��hH�S%���ۄ�&���K�0/���EVR�rSϓ� ��P��d�����7i��KT9v�0_ T�6�$֧�,Q�����?����~�L��i�����b��4�1�D5�l�|�q��i]�Q���Ϸ��\v��$>.UV�/�Lb�9����$9*Ѭ�ȝ;܏��Fb�I_	5����d��޳K|��� P�$�����.��r���猡{v�e�O�����>��*���ad<ʯ�|��c�PlXV9��g�F�v��Kq(��R(���ݝR(���ݡ@q+��^,8������or��콯��5sMI���f�+����خ�m�=���|vs�A����hɬ���>9t���R�^�G��2(b��z{Od�Y�E��n%�9��q8�� =�g��.�)��K�E��g�9�ƕi��g�_��H�l��/@�C�!�P��v/�IHM �x`H���v�����JE�Ơ?y����!���f����#�T:)�bQ/p��X_��<����]�b�m����� �Tg���L&D[^t�!e���2y�����8�t_H��&�ZBL��j5X�����D���J��-	�2����Ứ������2]���J�J�1�Y�X�Aw�|Ɩ�VY(f��ck3b�A��(lz��̓�\Zx^8�o
�)}ȴ� 3
һ�Z��l�I�,n�Gc�d�����Y��� ��S��24h�>��6$�ϳ�]rd�o�����Kq�L�P�"�,�!���ʙl`�H���?y�j��;��ϛ�aE�B�	����[L�[��w�.�7S� #��"b����R��T͚�D�Mp����ն2I $|}K�q�u�&�C� �����5�N!OZX�f~�+XƓ_]��(�hd�+�M�CX^�����|(ʁq��� rV��LOx��������D�von��R��_.������/���u.۰ ��K�-g+�ݤ+D���tp��T�؂Vrynz�j\�p� et���_�c��J��̴�,�WN�vk���Y %󣝜��i�H�H�	��Xhs���T��ȯ��yg��u���T$�X�i�hg[I6߾���q�Ne���G-��w�����<��/ �i�r�)�g�$G��?�KF�/���Z�Zs���V>�Ԏ�����oXI�NI3���yU�V�"ᒈQM�\�O�R6 �]��/C�������Z!�z�<�/6 @ݔ�
�4����!��$��.�zۛ����b����x��q���y���7��/+7������[������d/,N5�K,'\E�+���rjd����|����HI:p�:)�c��F]	��+�W8<-��%u5�
4�D�0�&%oe��׏ɋ�բ��[��!��K�W�����C��0\��kqIB�XK���/�)fL{/*��=R���h/��G�L�t�X��=�YKi�dn���dUF&ח(���ƫvp��kQ���%3u���_����Bx�K�U���O����C��''G�L��fg���#X���l��:���J��h��ؐ>��<�r�u�5W
��gĀ����`���X!s1�w������2C�`<t��z�dz�*q�
�h���92���}REe��>ἴ�&N���s���h9n`��b���d�������B4�e-7��?��7+�N����?��@MK_�h�Jʛ(�9V��	��?:b(�&��iq�-l�AW뫋���GϹ+ ��κ<3�	���tE�(���A���eZO՜��m�kcl�M�I�P���؉rW���|�����"#����V����=0��\��dz�ώ���b���?ŷ2�f�Teve�����a�%���`E;�n|6hJc�ɪk���-��!�ē��1�<0lrBg��ȉ� A�-�'F�!#�E/�o��/O���Q����7}!=@i�{���ak��V�핒����z����&��=�?�>�W�n��)qNO�~f�\JK�8�5)�Y~�b�� �h��]eR��]PS��f��m41�t@*u���_�h�R�X��]1�
W�=���xq܏�bi��SB��w����@����Q���dgo���ĘFH�� >k�#�-�c�2 c�}0�%,������
aة'��h���
V��\����q6U6p$���$���o������Nh�@+!LUN���d���N� ��4�1��NB.&�m����	/�u@u!�ku!���MEz:P�_�C���,Gd��,_3�`�f��*I��t��<b� XIcn��3P����4/�i����TQ�N�e6�4��K2�~�f0�ɠF�b4��D��W��� s���8�7�}{GT/��x���/��E}��ь�&a�1t@�Dh�ebg~J�@�/��k.���Y���͆VcG�¿�ȮVg���K�RG����aOG�yB�d,D�~Sd| -=U(�m�)D%�C����� n�J�%CG��O\)�h���%>,��L�
d�t[d�� ����V�#�K���4 �N�"���'c�ѫ���Y�轭�n�ƺ�Z�w����Ĵ��Hx]� >c,�43�T���b���ޛ�.nk��j���,|!xf�� ��L�+y`eg���]�o���h�G��[As	�~j�j8tܝ�Y�!�����n��a���)��+�_�[�&Ӧv��2����lN�����5/�կ�&�E&U�N{fy���6@��y�	�����	���'�����3��D�����'�M�I}���4���(�5Z�)E>?����e�������>�^z����T��M���c�C~rRz�,������S��\�,�
���!Ek
�Q���e)���,E������)�c�N�xL��c������%$"�k������#C͗��xnn����ʖ��8^,9�F���+��;| ��ܙ�i6�7�/^�'k'�'K���L�FL8�a�Wz����)��lA�J�~A��z������I�sO*����A�����[�"��ߕW�r�T+l}���l�#�M�S�9��F7�k�?@�'0PQO��5�j ����O��"�:{=.�����ȷxT�f^*rP��l��M�:O�*�7�*j�ag���b�DF	�����q&������%�h�^U��Ie �(�OO٫��C�y_���irq1s�5:@4���	-7n�p���?�Bx��_�89����,��f����:UMFS���i8p�J�����*��k��Ҷv@���o�=��ëL��R��DsJ�<��܏mo�z��L��{Z(B��'�l���В�NP��+�M}̔�17gV�o��'��MUR���/���׉u#��q~"���@�d2F���Ķ8�!�@�ww����04xj<,�*A�F��DD��?��,q�p	�Nq�־-cݠ�)\��Å&Ȱ�ɷ`���$�1����h!����-����RRND<�#Dc��Q0��'�2�͆��ʑ0��3��l˿��i�D�%��&r��L��B�_>o�.2j�->�}df���?��CAG���Շ
�`f�R��j	���)��AЊN��ֻ��.�U٭��ђa�p����H.�����Q�N�1�mX=��L�������bs: L��T]^pVb�.��6-��>��iǝI0q�x��
�5`%���Q���~�?ëֺ;�~���>CU8bф�@�1����E ��{:���P�͍��Ȩ�v|?����j�\��ŏ	a[I}=�������}�8���iյ�k�g�G�=�\�0�n�o�>�7d1h�� 7��u$)adYOw�,.�)t7�8��wRb�To��%�/lW��K�E�U;�[*�J5R�H��یVB�p{���i�w��~	�@q�B��gk��\X*2q6� ך;h�~�{�tU�X�*z��sD�h��\�w�O��ſ�T\l$���xp���7�DM�v`�prc�@+d
_�ʮTw�X9�����AG#D��]f��r��a��S�Z��}h��b�R珘�I���T�����z.o�p����K���ȌxVj3��\+h����i�CfKcKYZ�����V�Eׯ��~\�M�|�
J-�M�!�0(���5;X!S��������G��U�� �Dkp������j4�P�4\�"�Ӈ�������V�/�xFCv���ϠwZMI25 �{�O?��n3���V���I���"k]�%���a-a���*���c�@�j�{���5T�3)<P|n��rN�$���hj(��Fx���/�����QLKN�V���v���( @N�}���ӳ	n���lB���R��	���|o tD��6�0y�ż�*���d����O���q�h,���4d�EeF��6SsRs�%A �|Ӱ���j��#�M<Z#.��\�{��Z�2���$h����De��+�����C-ѭϩ\T��w{�|0�P�$(h7P8nt���33��%�c�zOv	�q_>^�>lo[�K��n�YH�+�����%Ի�X��7h�;���ne4��FJ��yz�$U%el��_>��@�\������b�5��&�����ԍ}ږ����lҜo��݊V�u��-��9qi���3�<�����G�U��4����R*��ځ����O	F���m�+����t$�,��A3��tl�����=���Z}�V��?�����X�?
� ��j1�uD���x�HZ��}(ww�������#Ij��&	��3ZMK�Wϊ�#r�|�~N{�1(�(jq�91J���z��U΍�~��z[:��]�]�w����9�<[�Zh�E��l�.��i;�u�GgAՕ�"�['΋��lC	-����I��s*I7o��2M�?�%2}��Ӱ��<��S[�?�>#X�6i�A '�"�ez2T����]j�;�hc�����-��ֳ���ID�z��a�T��O��|�|�e�Q	��ᴃ�v؏�L���@�u��o�Y%x�D9.��V�1�3�~y���y�+�6���ַ��CpZ�0�u�`P����ʞ�X	��q?�P���'���E�y�٥H�G�R�a\ϫ��P��:�8��m�G;k���vXs:�mk� �&��]�Z��R��7�`����%�>�MȐ����=�`N?U��*����I�4Ո	K;���x*�9��M������8�4���|�⬽�!����;�6��𛙴����5('0�p�7�����ͨ�o�i���Ӿ|-ު.(D�Ր�v���a<��ڄUU]��X?����Z�y���k{�StȌE��6�:���E�x���$�盄��Lt��5�.Fㆆ/����')"��zOY��x�C�������n��٩ɸ7�$6��q��#�I�M63�oe��(Լ<T��yjR�G����VG�ZrB"�����?�>g痏��9���P��^FXU+�P�H��K�/<���l!~TM�"X�t���T=����W������K_$��CiBn+-�j�LC��s[���.�[FIY�|ʾ�YJ~~XA�ο'~���e�r=�e���_��RiCM�PR��Y"��D0y�]�CZ��l��L+4���ML�!9�T� ��S��c��h��-�#�]���ppN�����M�V�`�4�^F����-̓��Y�X�������j����B@JV.O�밋��������K�7"j�^�ʒ���I��bHH���BFa4�[��D�����A���Z��^���!ÿ�I�Q���`���������Kj֛�釄veD���[�� e�9ՅI�~j��:�p=��]����c����6n4�ъ�k[��|q��i�6��,��^��f���>�x;I�ը��5Q����-<���_������^�*��y'b����6�o}6��2����6L>\��&s&��<�c����¡�� �E�t����n8�bd��7I��M^V��α..�3J�:�li�mz۰�͵�X�7�o�#
S������@�n%`3��^�~tvQ�`n^F^ZBZn�&D�������/�涽D@`X��O+)EE��1i��N���T۬�I��G���X���fT�|���M�%�د�����X����ѱ2�7!7M�Mf�7��/qM��DN)�ti���ū!����?*A� ��U������B��{�n��{K�/\(ưˀl����;�`�`��:?|��3�������|�7ДT��[ ��nǈ��7w�M#�%�dY�p~�}�F ~o'u�S�稟��3K�e����q�pk���'r�Μ`Ѧ�f��� �
�k.6��g�;}��8E��]b�v��{~ ��fӷ�YX9\�E�M�B��c��pL��!���X�����!�p���!�[%y6Z��^���W�)�g)b����_�S��jO��C�iK�M�ֻb����*�К�3�sh8/�Q^�谰ܫ�����du�A���d?��hf}�Y��sofj[��k�}�b`������f��'��m�������a!W�^lĤI�6���z�'Nf����t��/4@4���ǰ�!Z��KRR�̿~ܞ��EP�AߔSb|�{�G�"A���]|U��or�qPb#u1���q�o�%"]fl�`����^�wmZ�Bd8��A�Q��M&�r�P��R� ���؂c)�Z<%����+m�\خ�?;3#��3Ѷd؊�8��f<KdM#�WYm�_(E�%�LKqg�ۃ�`�[�o���,NtI�J!.Y]r�A\f��ǳ8�[0Gf�W��#�I�gS�6�룮L!�Aq��z���[�o�	"�׳�ed��.�)��^��F��c�.�ö)8X��,v��I�9\NH@{Pd�z���+2�"\Ֆ��{G�P��?����'�9)`
��T$��5����6�0.���G��m<��w�z%�:�����2ӫoL7��E,_zl�p����� �Q��a�9<��6�I��&xx���j�;۰K(:<���k(;��H�����3�����ʛ���*��^����ͳ����k<ߪ����"�I��|תR�(����?���TḚխ�lwB��N��47�T��@�5gSp/>�<�e�n�?t8��K��[x��K���ƹ�j�>��:�i�4��^E��WT�{�)�f�X� 2s+4���Ѫ�qZx��)�Bo�����U��-��Ǳ֤�g�^����<��#5�2&7�-�౞! �F��X����d�	�/�J�B�&�N�e^��D5vz��ӿo�i�
n�In��v(�*�=����4B)�a������G�k|5��=&ϳ�6�5M�ӳ�-ɈF�G�x�7�L�S��yR@���/��Ȫ��F�nL��?v��q_ wbx���4 ��d�c}�7�~�z#�B�O%��[�z47�B����5͜���R�ZLN!��h-�,�YB���o�#�%ܱ�/�a����;Z(���beS�6�h������mv?��@���Yn���\MY�?�K� ����Г.p,�d�9�Y KG���zm�_�lu��|`A��@0�w���%`�Y�S��' ��S�L�QJ�%�y'�^���&y�������K�難6g/�Xb���9uai���NE��O�- �(�9��!�a�w���>������6Z,����e~�{�~��ï)�ýZ2����Ż���)��A��ck�ٗ�KcE�ݪ9�o���?֮J�MB]9\ƣƹ����lT���s�|P��{�J3��������T"����P|����F7Ag���n�5�g�~��ƹ��q��x8Uᭊu̻��Ċ�o�WS��.Ud��|�ɝ��\�OÎ��K7��&&v���X�W��G���$<���C�v! &���~q�M�&�btNJ����>�E�Ŗ�V�t��57�"�q��˧�����F�B.��w�������n7�S�B�ܗ�"�!�4:�e�Q=O5�[�-����H���ϗ뻶߱�d�-�Mq���oTS-p�p�BF���&W�)�hT��0§&B�}���X�ege7Y�����Tc�\������}F�BfM�g�����]�]�[�>����?��|I 6�����M�t�X�w���е�0[����x��h�����VƱ�YwqS,W~W{a$<�t��~d�[Z�"���x����˼E���}l*���y4$�z��O�.N�iW`C�7q�;XL������ʮ�5��B�-D��o򤞯����͚u:}[8[xz^G�C1�G��\���Ƴ����8}s��*Ͱ��@egcr��P�֭���M��K�� ��B�^f��nǱ�K�t��W���_ t,S��� �a�fC�v���D�BG�PV)����P_\�6l�_'�~�,h�Y;��IS逬G��	�=�� e���X��g�c�js�nɦ!��[�(4����a�h^X�q����]�Q�.þ(<�{i8���kO�֡fbR�ZY�"*��P{�?xy�֜K�T�*�ŋ��l���Q�E���Ԭ�kXՒ�(O��"1Fm�IF��G<�d�-Wy��;3	�{Tи����'G&����Iؼgn$v��YC����l�{�����Ҿ�z��Kg�R��>�W��W���mt�34�s�������d�H,b�z�z����5��<�z����)呠?�ː�LZ�|<�LJ� H�(Ns|,F6��iz�<9F���q�j�\�M���y��>�Ҫr����<�b��X��J�)��aK)���Lű(򖞉�4I�����#:+�%͊��wk�qO��Ǭ�V��hZB�l}�����ub�������7da�yMvM=E��õa��Q3&�(m�^�+��iv��%�`|7��*bw򒢢9F�!�}}���Q�zDlZ�?�pR\W�C� $�q�O�?���~a���w��'D\TǨX.�8I!�~�M���i����8���׹]J��B6#������W\�d/
t��5q�V�C"x�S�2`� mo��-8����v�v�nr�
Y�S[��Yr���E�Y�$�C2�R�@SF�L�L����Ŷ��g_�i��J��\�<ެ�G/yi��\�-�E�{k���ײ%>��ЄR��2�{R]����+���3x��!���gh�6���O�p������E�ħ1\y��)=�32?�����Q�k�9�X-a�''���j!/F�G�jF�/��N�j�sP͑�<L�|����q2L�r��g�S�9�e)�~����6�oG�B2�T6~tTR˗1TE�k��d��!����).�?]8ƨ e�
�����4	a�By�7U+�KEC5BE�N��*�`�(���t-���xdEG�F��/;��^u��ԓ�"�[�s%�"�  }Nu�N9rfա��M��l�"�m��NvOː٥��b���o��}2I@�N S��0vۻ�J���bӑ��ϛG$km�D�M��aӖ;m+��bh�A�7�χS�]����={{�Jq���DX,�}�v��ͱ����<�jj|���_D 7/%QB,'wJص�W����{���a �*�8V���"+	�lA��)J[Y��i����n?��"���6a�V��pǉ��(%u�	��(]-����n�+��_R,��o�B��.Г�%��uHw6�ܙa��/�x�j��X��E��窋�����㭯�FC�I�y��A�.M���tc�S��w �P�S��׏����+���n>s�Z���\M8D�S��t�DEL��܏��oܞ�ӳ�	>w	�����n������*���&l�J�>������I�<Y�E�D~Ôy�����֍�3x9����iaa��E��O<�?�/��X8CF�e��]U�&����gɗ�Fa���zy��i�c�?N�<A3i@5�ߕ��l]Ei�+x��-
m��=p"C1eA4Yg��w��KY�˲^�ym
Oh�%�ٛ8�� �0�Ts���m��`�Ul���԰Qi`���?c��yVL�D ߲h�C]g]�/X��@��ֈ�Q�L��38 Ī�k��ބ.�>ǣ*Ju��6����#��Dc�rz�l(v��!F۪?��x�~�SN�T3�� ̘LmXo�Y������i��DA�_2w���/���_U% h��y2a�N��(U#%�~����Hl-R8ء�K��~���tw�C�p)ϰ��/����訕�s�
�ZՋڥ �C�e�� ����HK���K�4�+t�d�5�H��t��;0JX_=�:������KH9�2Ś�쇀P��h��7Q���x(�a���p���(3?1F9w�)骤&:�/��_�kX�g��3u�?�5Ag͊�����M�_��BðѼ�k�>�������. P��UUl_����s���t�L)�׹�D�8f�w���b�ܚk�H��>}sZ��������]7o/��c�) Jj%�����y���$~�Z�CI��Y3�nj�>�_JnqQu�U�|7��A�&/Z��XFY)���6+�''��q����DB��T�:�����6h-�Z���ס�U#�13�$�;��*�RR315��͛l:�r�Te�t#�I���ǣ��(�M�I'�8�g��$����W�J�>�_?��#u�ݤ�jhr�}~K,l�*6�Z�^��'2'�Kd�]�.��O���HҞ��\���a���na�ޏ�������~B� ņ����V��wU�V����a��5�^��Ck?i�ı�� �k�'�h�p\n��Q��,!.�bc9�8N�}63�;V5Ϙz�[JU�s�G���.1ʹ�����GX���DXYA�<A�xx\Tm��7d�H�E��h���78
�	ˋ��kܦ�!8��/l�c���o�(�@%���v��������<�����_���ڍ���^"n.�+uZar�)���{t~a�f'%r���@ ��&�h��"� ����^��Tc&���c�@d}��NH)��qh�Ymw/��H[mYM9������L�Nژ���5Yc�� �Ҍ}٘쭤��31��F�equ��w*:��m\=`��(r]���E�q��r�A>�fq��4v�z3�}G�̊�j� �TVy�7�]���)�0��\�a.����ČF�)ғˬ�Е@wNm��MR�I����J������bRrVn�p�E�.���aIwR�g|Xqw�fU���5jЮ���t���J���U9�P;A;嘔_���X�bR�o��}��æ��u�5�L�ާ��%�����Ϟa�[8��! ڹ���/Od!����
do��0��J�;;�u�﫶ϐȿ�#��7��(�
K�L�'�CY��j�xw�W�[��9'(qJ�� 1Q���_170ٲ�ao5~����^�3�2�EI�@�~4���f/FK/�%�IV�E/%7{�����)�.���3%�鬤uu��(��3�������ѯ��>�k��#S�tF\�6���v�����1�`��t]]��@x��?h��=��t$��B�8�خP�۷�K�N*	��`�ޢ�H�;�z�"��=���_�mh�-���&�e? ��>��7�'玫�Up� b!bh��#@�ocw9"ng��g�8�0����,n�ވ�7y`�ݴ����n�xN�� �S�Ԭ N���SƓ����Y��ȧ_��rmb##��3�.�6V� d-Q̍���Y�����><��_�5���
������dȢ�J�_�.ܦH����m���>g
�����]��=Ŋ��^7V���E��SQ���F���]k��������C�v\k�+}����@|\s	t�?���R��+���ϸ��8W�t����+-�sB}iHl�V
Q�KzU���n�5�%���T�z6wV��멫�Kv�-���{5��]N��w��� ��?��x�Y"�Ll�]�j�H9
�%z������O�haE�Lӫ��F�ͯ��e�x�+:��I#�?�ظpq��:�#�]���������{���o&{xH"���֑�3�Z��u	E|*B �W����4ڈ3�����o]C=S&��_AȠY�un����O���<LD9�oE�_���]�O*:�EHt��9���a��Ej)��k*|��P���_@�i��|�Ҋ�<!y�d�Pv�T{=�~��08j8,�c�@���#��KgS���Ϫ��c�Bo8n��^Q�'�y]�E�p�*�7�+{���e��3�<_��$�f]�1Ą�����$7?{�lg۶�o�^Z�����LeI�6k=p��2����6�m�n#�[����_
���r�_}�+ժk�{��Pp�7��Q�b���5��gGd��@$e��C����s��wk�.��S�R�"7�����fE'�e��I:� '�<�����C�4l4tTV��pO�y�5:��b���C�C/���o�o���`x��U�i��l��m`�|�܌
�Hq{���-�A���R�*��L��Z�*��e^C	�y`e�9��j�����Wrl�%�?i�`
Q���!X���p`�2HPbo�ɾ= zt�#hШ�jVb#�g�d ���J�N��uk��B�1Y�6k nre닚�鮗��ӊ7jپ�輭͛5l�1J�Y�i�1����J`�s�:k�5ص_������P�!95��-���^L
�/1D���d�������k��|�~���v�]13�2�����
�^q?T�#Xܽy�ޢ�D�F9N�yż���n��ʒ��v
����<�)���}��Q'��,�<��Jž�����J��˸+���=�?侬e��)�I�e-e|>dv��,����)R�:����O2��k��}DG�Җ�'���(^��=)2b���٦|J��/_ˇk夨I��$�#���\H���H*�=��q7��*��yʧ��/I~�߯����G��^\@�A��-�ET;��9�0�D���w~l��l+�c�)\M\�@���E\V�g>}uf�Y��$7��p��2J�Հm/�Ɛ��`��e�^�b���_Й�P���ҫi��D�^N��z�}�Fp\���e��64>�4,�'x�T��l�����T/� ���br����όE�;�(�;6�s�������mm���Ѯ�D�m�Z��l��y�FAG>�^���P�V��-\�?g<*l���(�-vl�����+o����Q:8d6>��^n�������s,.�d l�oT�T�y��`��Z�/��B�J�՘�/�8Ӄm��m�\��#���R�N�W�:m���|��M��j���s�I�$�����V���d�X���@[�ϴ���}0}C?A�'����b"6/�i10L��;<�I��0.����6�^Hc���%���	��Z�C�I����g���8p8XR
M�o�Ϛ)�gi��'^/r7�=�hJ���<|\:R�6>�iQBaz�ܛ�u���z�Q�(�e��iRD;Y �Nn�C�=/�X<^6 �r��I��4�W�_`�v�z�����3N[Չ���}� �m�­�w�P��5t�����TCΏ�
K��]��E�`�����xcAط߮z����N=�~���y���a^@����LH��6B ��ϦO����y�i�s��[��3��AoL�H�к8�&24�2P�1�Yc�;�s-���3�"|�;'@C
��g��Q�L����'sl���&w�3�S���� PK�ZV���!�c�d'σ��6��3����2����e�K7O�JF���w� ���%Sˡ~�������2w�4$=�ƻ�Fa'���pE���u�dX�h���2��L�tI=L���������y(��l�-سr{N��jr��7
�G�*��K�2���A��T�>��a�ң#r��>�1�ԛ�ya�X瑫�'��4�����j��^����0���$�mV�ȇ��$R�&��n�Z�;ߺ�V��h�舡�/_����N �_�Q9���:tֲ�7Q�S���2�R�v�w��y(=�뜯��9�ǫ�!X���`'�@�����l�j4q�j�DP�������+�bq����IR��ne�O���pq��<���9�iU�}2���d��`��"���Į���翐L�����Q�8SEj�|�̦��V�ݭ�&�o�����ﺪ��������3�h)�w'��a/J44�(k�f�i����t�<EBQ=�?��*���+!b��v�n���ܩY��ԏ�@��Z�*���L��L������I>6%�R�;�!��$�ߠ�z.�1_���!sԳ��ϟl���+���R(�0�l5���'�y�%�5[L�*6�]ַ���;�a[^31�����8����4?nf_�['�J�Ə�R�-q?NbE�9�2���� ��(\=q��2W��.1�H�M���Ԭ2�A���&��Ҽ�k��*�;�0|���d �u��I;��x��RO�h)d��A���o�[�jp�{�G��JD����Q�'uL:�?Ʋߟ)�%1Ÿ�W��C"x̩-�:L�C�{i��s=�,^_k��* �TB}��<�WC�w��Fb����u�+ps�?� ���Z�K���j/���A�|(�)ð\:�)��{�z{�ݿ�R�Q�-��$8E���3�2Z^��6�&l�5�gS�R[Ӻ�)��6˿g	d��Zyk�C�o0�vㆀ%)v�)[�d����t�w�t?���		�+H2b_Ք�m:�o��`q�a=CU�PtL�����k���S5؟r\���ر��Ez�D��p�����r���}Cy)SS��bE����ec����e�F���A~nf�~���EX6�TA��]�w��Y#�c���los��o���}p������/���ce�@���d�bc��#�F���jg`���'��*tlmgo�>��Q5W�n8E�KLo�gq�:OOCӞ�[;׾$�Bh�[#y����UZ�^��@��.�&�TKLI�j�3���.��Fy��I�^�	|�r��4ƃ2��X8X8��=��?hty����b��=��ڄ-Zݠ�'J*�|�u����*u�°���mɊEN/I%��ny(����� ̘�TE9y���������Σ��d�&��:%��⋨��؋Kp����El3,��.P=�za�]��׀K&u�R���%37�Ĺ@)^'_���?}L�:�<6�+������4����X�aŇ�}�/K�BJ��A0��9ͦ�;O��]�t*[�
	5�W;�圌���M���{.;�h������@}����s6dh��k�ǉ���7���)�`w���c�hdD�R�tm�m�T������V�z8�{-���n�^����5E'G������I��&�'��o��I��nz�1�/���"C�G�\6T��n�_������~����;~��'hb�;o���k�ۄ�i$�5�gX��6$K��*K,����9H�L��V�TI,3zi^���|�T�ˌ�}Ԣ�>�My谉�˭E��c�v*��\s�ʵ�m��7��c �u�\���X>��:�'�c1�b���7Q�s�8��"$B9�`�����/� �&ϊ+L��G#�Dݶ�%ᙦ$��K��7ږ0?"�ӟ;�w�⽸JIG,�Mi�C+�4:=�c�S6�`q�ġ�B����$��7���kF�Dq*u��AS���a��*n��x��Z+S~�w�|�%K��D3@��>��p��z.��:14��A��vjz����e�<kl���  �sc}��_���d��� H���X�m9@�濫�����H�I����!��
a\Jy)TN���3O5���ZF�A���꧑P�����y66ܛP6���U4���"��q�p�Z�w�"Kh'�7p�&��.
��\����Ӝ�]���ye��j%k]���R�l4��yHz��^��.�.\Ez��$=ME(��S�t�"�=f��ݡ¸�����<���	[��>W��KD��eT
E����hd+��h�Jo���rieo��=�ǝ���JqmK@����١�g�i���*y�����R�����y9�C��(8VT�cm��ypHo����VnQ�e���m@�b/MM��0[~]?#����:Xx2ڳ�&m�&0)�����Ͽ�m�s��{.a��Æ0�|�'�0��˒1̳�4� /�����k_b>F���2�\�7�����E'N;��zt �Q�&�PQ�հ�ȆH_�^�Ðo3�����U����f&��p�+'+��ރg�s�s�$�E���~�lF���Jm-J�2eѠUh�L��R����ϡ���0�l�V��9�@�Z�S&��+�!lh"ǀe�ˋk��{}x��R���p��r/fX���b��=41i��4������0�٦�=�^��ȶ��yE���d�g|`�/�p��c�`!��X7���}5.�!��l��~LtNx)++?W�I�ɲ��~���.v�"\����m��䗮d�j�9Dq��}X,x@L�/;�8jdX�_��3{�p���r��u��?�~R��,�h�*[ÖT��R� Nc�}�ݩU�
v��������Ġ�>g�}�e`�m~��a�/�+�Z��T��oT�!�]��/!D�ך�ǖh�������~���u'�O`e%��X�릠AGu��`���Odsf}ƿ����:l��ۈ���-�kml��zO���!5���G�E���#8V��h��N�S�ܥs��kW��wJ�5�>�!��?��Xm�iz��g�|���u�3�Iц�CǾ=��~?V�ܱ���嚣5���+���ȞY}%���{��������g����|ߑ/��f��Zm0��ܻ3F2lN<��8nN(P�,u�G�=��Ĥ���Y���h4������/��QLM���n���:��Gv�N�^��%E:��5�b�!#ʲfB `�?a?e*��`|!_�Wuw�ݝ�#����B���փ������4k�l+Bf�Y��Ðk���j��}��1��	L������v��c��H�7�eEez���0��Μ"�����?����[�[������p@Ď(��=��_���/>��Y听b�/��rp�,�P5����F��V>�p��f�l�APTEQ�!��k_k�m���&(гϾ��WmͶ'��DeyeRb0AŪ��}C}����n�;���EM*,�뿭G�UwT%�lͶ���x�� �`�;�r�3���  ,�i��D�d2��㎧}z�b)稳zO���� ��b��su��%-�-�y�Y&}�aps��/���[�Ϝq���zC�޳����������޹o����'v�����_��XRP���G+�+_���7��,v��i�$Byay�_k׭^7�rB���G�߽o�W�N��h7��PuG�]�wut�5��_�!�|�]�EL�i���y9y���+�V4v6���X��.���"Z���m(3��������ƞF X��à��G PF�'��PQT��p6凩/z<ucB@q���m*ؤ�a�C�Xm�j~埯Hxr�!�k���bo�k��Sq��ȑ@(�y������3b�H�п�O�1�5����{���k�פ&�Z�3�@��}���|��Dh���yCގ��c_�9�+�DQ ��Q�����ͩI�Sc�щ�w�����{dڽ(�ް�o�������u�7G�x9�(   ��ǝg�p����,˓�3�{D6�/����ޡ���Ρ�!M�&����ƀ�+���:y�y<��8.h�/ ��G�&Ѵ:kurbr�:��a��8z�V�v���"��r4(%,�U�B(�<�;Ի)S�%Q�Ш/n��y�ߣ�׋yE�R��=xa0"Er2r�(����v��[󯚋��0��������W-&�3�IIL���1��&��Pr���b��������QJeUI!	K�^oL�����84�)X�T�0���#��xQ�TESd,F��h��]��x �q��`"���֞�-�d�"sq��7�}�ͧ�l�R��W�/�&��؅��.};<Y�[�[ު}���}�&g0��1gә��9������eT#��ȧ�O�X�b����Ό���s9 AX7w7��9�������p9�}�oׁ]ޠw֢u���峴�~�u�2�x��q�(����߶�۶�n�5ٚdIZH�2����v�>��d�ɨ�+�4� $�	f�� 0�%���T��AȚ`�����~uߖ�-�V�ӷyEQ﫮����f����������r��30�ds�E�J�j4�.�7�L(TU�@��8�["��1ۚ]����;��eU�5=9!�b��l2���9�����c���8[�Y�R҇����
����KJJbJ�5�$�
r
�rc���JQo�;�`�M&���~9tJr����@��8�[b����������l�rk�y�y�6�Mf�#�i��J�Q���^g�������~RصH@,F��=���k3h��R�qܲB �ќ��_�[�*k�A0`�9���&� �C���E����7��8���0&i�=8<2l2��E[
QTU�����&�8n><��8�����1�`E�ʵ?�����8�����Z~�qK���q�q�-�� �X��4�;    IEND�B`�PK   R��T1b�!�  �     jsons/user_defined.json���n�0E��Z"D�aһ �d�"H�Uaz�)�TI)�a��;��E�@�� Ν������FK4F~��X�[��'��
.0��8�I������ڤ^�@�T�~�a�h�Vi��d�ʚ2��B4g^�5g�j�ҒjU�IN���!����+�`��`����63�w���[w�G�r�fec�U�[����X	E�N���jň:���=�w�~�<�,	|���g���B�s&2"K�(� ���5�|���E���I���y4�F3:�6U��i���=�M�c�$�tz�s�����~����x�pG��:�e��.7�]�q����B��a�Ü�0��V�67�"9+M�KS��PQ(b�D_�9�9�!�.ȹ�p�-�ˣ����"����������9�9�~&<���g��
�;49�n���PK
   R��T�FT�G  �)                   cirkitFile.jsonPK
   Ǵ�T��v�({  �  /             t  images/44c8d6ed-f4a1-42f0-8f26-136091f6581e.pngPK
   '��T~D'�K #L /             �  images/838b34ec-6803-475a-b54a-babfd323e900.pngPK
   R��T1b�!�  �               � jsons/user_defined.jsonPK      <  ��   